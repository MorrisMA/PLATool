`timescale 1ns / 1ps

module PLA(
    input  Rst,
    input  Clk,
    input  CE,
    input  [8:0] A,
    output reg [35:0] Q
);

wire    [511:0] P;

assign P[  0] = ~A[0] & ~A[1] & ~A[2] & ~A[3] & ~A[4] & ~A[5] & ~A[6] & 
                ~A[7] & ~A[8];
assign P[  1] =  A[0] & ~A[1] & ~A[2] & ~A[3] & ~A[4] & ~A[5] & ~A[6] & 
                ~A[7] & ~A[8];
assign P[  2] = ~A[0] &  A[1] & ~A[2] & ~A[3] & ~A[4] & ~A[5] & ~A[6] & 
                ~A[7] & ~A[8];
assign P[  3] =  A[0] &  A[1] & ~A[2] & ~A[3] & ~A[4] & ~A[5] & ~A[6] & 
                ~A[7] & ~A[8];
assign P[  4] = ~A[0] & ~A[1] &  A[2] & ~A[3] & ~A[4] & ~A[5] & ~A[6] & 
                ~A[7] & ~A[8];
assign P[  5] =  A[0] & ~A[1] &  A[2] & ~A[3] & ~A[4] & ~A[5] & ~A[6] & 
                ~A[7] & ~A[8];
assign P[  6] = ~A[0] &  A[1] &  A[2] & ~A[3] & ~A[4] & ~A[5] & ~A[6] & 
                ~A[7] & ~A[8];
assign P[  7] =  A[0] &  A[1] &  A[2] & ~A[3] & ~A[4] & ~A[5] & ~A[6] & 
                ~A[7] & ~A[8];
assign P[  8] = ~A[0] & ~A[1] & ~A[2] &  A[3] & ~A[4] & ~A[5] & ~A[6] & 
                ~A[7] & ~A[8];
assign P[  9] =  A[0] & ~A[1] & ~A[2] &  A[3] & ~A[4] & ~A[5] & ~A[6] & 
                ~A[7] & ~A[8];
assign P[ 10] = ~A[0] &  A[1] & ~A[2] &  A[3] & ~A[4] & ~A[5] & ~A[6] & 
                ~A[7] & ~A[8];
assign P[ 11] =  A[0] &  A[1] & ~A[2] &  A[3] & ~A[4] & ~A[5] & ~A[6] & 
                ~A[7] & ~A[8];
assign P[ 12] = ~A[0] & ~A[1] &  A[2] &  A[3] & ~A[4] & ~A[5] & ~A[6] & 
                ~A[7] & ~A[8];
assign P[ 13] =  A[0] & ~A[1] &  A[2] &  A[3] & ~A[4] & ~A[5] & ~A[6] & 
                ~A[7] & ~A[8];
assign P[ 14] = ~A[0] &  A[1] &  A[2] &  A[3] & ~A[4] & ~A[5] & ~A[6] & 
                ~A[7] & ~A[8];
assign P[ 15] =  A[0] &  A[1] &  A[2] &  A[3] & ~A[4] & ~A[5] & ~A[6] & 
                ~A[7] & ~A[8];
assign P[ 16] = ~A[0] & ~A[1] & ~A[2] & ~A[3] &  A[4] & ~A[5] & ~A[6] & 
                ~A[7] & ~A[8];
assign P[ 17] =  A[0] & ~A[1] & ~A[2] & ~A[3] &  A[4] & ~A[5] & ~A[6] & 
                ~A[7] & ~A[8];
assign P[ 18] = ~A[0] &  A[1] & ~A[2] & ~A[3] &  A[4] & ~A[5] & ~A[6] & 
                ~A[7] & ~A[8];
assign P[ 19] =  A[0] &  A[1] & ~A[2] & ~A[3] &  A[4] & ~A[5] & ~A[6] & 
                ~A[7] & ~A[8];
assign P[ 20] = ~A[0] & ~A[1] &  A[2] & ~A[3] &  A[4] & ~A[5] & ~A[6] & 
                ~A[7] & ~A[8];
assign P[ 21] =  A[0] & ~A[1] &  A[2] & ~A[3] &  A[4] & ~A[5] & ~A[6] & 
                ~A[7] & ~A[8];
assign P[ 22] = ~A[0] &  A[1] &  A[2] & ~A[3] &  A[4] & ~A[5] & ~A[6] & 
                ~A[7] & ~A[8];
assign P[ 23] =  A[0] &  A[1] &  A[2] & ~A[3] &  A[4] & ~A[5] & ~A[6] & 
                ~A[7] & ~A[8];
assign P[ 24] = ~A[0] & ~A[1] & ~A[2] &  A[3] &  A[4] & ~A[5] & ~A[6] & 
                ~A[7] & ~A[8];
assign P[ 25] =  A[0] & ~A[1] & ~A[2] &  A[3] &  A[4] & ~A[5] & ~A[6] & 
                ~A[7] & ~A[8];
assign P[ 26] = ~A[0] &  A[1] & ~A[2] &  A[3] &  A[4] & ~A[5] & ~A[6] & 
                ~A[7] & ~A[8];
assign P[ 27] =  A[0] &  A[1] & ~A[2] &  A[3] &  A[4] & ~A[5] & ~A[6] & 
                ~A[7] & ~A[8];
assign P[ 28] = ~A[0] & ~A[1] &  A[2] &  A[3] &  A[4] & ~A[5] & ~A[6] & 
                ~A[7] & ~A[8];
assign P[ 29] =  A[0] & ~A[1] &  A[2] &  A[3] &  A[4] & ~A[5] & ~A[6] & 
                ~A[7] & ~A[8];
assign P[ 30] = ~A[0] &  A[1] &  A[2] &  A[3] &  A[4] & ~A[5] & ~A[6] & 
                ~A[7] & ~A[8];
assign P[ 31] =  A[0] &  A[1] &  A[2] &  A[3] &  A[4] & ~A[5] & ~A[6] & 
                ~A[7] & ~A[8];
assign P[ 32] = ~A[0] & ~A[1] & ~A[2] & ~A[3] & ~A[4] &  A[5] & ~A[6] & 
                ~A[7] & ~A[8];
assign P[ 33] =  A[0] & ~A[1] & ~A[2] & ~A[3] & ~A[4] &  A[5] & ~A[6] & 
                ~A[7] & ~A[8];
assign P[ 34] = ~A[0] &  A[1] & ~A[2] & ~A[3] & ~A[4] &  A[5] & ~A[6] & 
                ~A[7] & ~A[8];
assign P[ 35] =  A[0] &  A[1] & ~A[2] & ~A[3] & ~A[4] &  A[5] & ~A[6] & 
                ~A[7] & ~A[8];
assign P[ 36] = ~A[0] & ~A[1] &  A[2] & ~A[3] & ~A[4] &  A[5] & ~A[6] & 
                ~A[7] & ~A[8];
assign P[ 37] =  A[0] & ~A[1] &  A[2] & ~A[3] & ~A[4] &  A[5] & ~A[6] & 
                ~A[7] & ~A[8];
assign P[ 38] = ~A[0] &  A[1] &  A[2] & ~A[3] & ~A[4] &  A[5] & ~A[6] & 
                ~A[7] & ~A[8];
assign P[ 39] =  A[0] &  A[1] &  A[2] & ~A[3] & ~A[4] &  A[5] & ~A[6] & 
                ~A[7] & ~A[8];
assign P[ 40] = ~A[0] & ~A[1] & ~A[2] &  A[3] & ~A[4] &  A[5] & ~A[6] & 
                ~A[7] & ~A[8];
assign P[ 41] =  A[0] & ~A[1] & ~A[2] &  A[3] & ~A[4] &  A[5] & ~A[6] & 
                ~A[7] & ~A[8];
assign P[ 42] = ~A[0] &  A[1] & ~A[2] &  A[3] & ~A[4] &  A[5] & ~A[6] & 
                ~A[7] & ~A[8];
assign P[ 43] =  A[0] &  A[1] & ~A[2] &  A[3] & ~A[4] &  A[5] & ~A[6] & 
                ~A[7] & ~A[8];
assign P[ 44] = ~A[0] & ~A[1] &  A[2] &  A[3] & ~A[4] &  A[5] & ~A[6] & 
                ~A[7] & ~A[8];
assign P[ 45] =  A[0] & ~A[1] &  A[2] &  A[3] & ~A[4] &  A[5] & ~A[6] & 
                ~A[7] & ~A[8];
assign P[ 46] = ~A[0] &  A[1] &  A[2] &  A[3] & ~A[4] &  A[5] & ~A[6] & 
                ~A[7] & ~A[8];
assign P[ 47] =  A[0] &  A[1] &  A[2] &  A[3] & ~A[4] &  A[5] & ~A[6] & 
                ~A[7] & ~A[8];
assign P[ 48] = ~A[0] & ~A[1] & ~A[2] & ~A[3] &  A[4] &  A[5] & ~A[6] & 
                ~A[7] & ~A[8];
assign P[ 49] =  A[0] & ~A[1] & ~A[2] & ~A[3] &  A[4] &  A[5] & ~A[6] & 
                ~A[7] & ~A[8];
assign P[ 50] = ~A[0] &  A[1] & ~A[2] & ~A[3] &  A[4] &  A[5] & ~A[6] & 
                ~A[7] & ~A[8];
assign P[ 51] =  A[0] &  A[1] & ~A[2] & ~A[3] &  A[4] &  A[5] & ~A[6] & 
                ~A[7] & ~A[8];
assign P[ 52] = ~A[0] & ~A[1] &  A[2] & ~A[3] &  A[4] &  A[5] & ~A[6] & 
                ~A[7] & ~A[8];
assign P[ 53] =  A[0] & ~A[1] &  A[2] & ~A[3] &  A[4] &  A[5] & ~A[6] & 
                ~A[7] & ~A[8];
assign P[ 54] = ~A[0] &  A[1] &  A[2] & ~A[3] &  A[4] &  A[5] & ~A[6] & 
                ~A[7] & ~A[8];
assign P[ 55] =  A[0] &  A[1] &  A[2] & ~A[3] &  A[4] &  A[5] & ~A[6] & 
                ~A[7] & ~A[8];
assign P[ 56] = ~A[0] & ~A[1] & ~A[2] &  A[3] &  A[4] &  A[5] & ~A[6] & 
                ~A[7] & ~A[8];
assign P[ 57] =  A[0] & ~A[1] & ~A[2] &  A[3] &  A[4] &  A[5] & ~A[6] & 
                ~A[7] & ~A[8];
assign P[ 58] = ~A[0] &  A[1] & ~A[2] &  A[3] &  A[4] &  A[5] & ~A[6] & 
                ~A[7] & ~A[8];
assign P[ 59] =  A[0] &  A[1] & ~A[2] &  A[3] &  A[4] &  A[5] & ~A[6] & 
                ~A[7] & ~A[8];
assign P[ 60] = ~A[0] & ~A[1] &  A[2] &  A[3] &  A[4] &  A[5] & ~A[6] & 
                ~A[7] & ~A[8];
assign P[ 61] =  A[0] & ~A[1] &  A[2] &  A[3] &  A[4] &  A[5] & ~A[6] & 
                ~A[7] & ~A[8];
assign P[ 62] = ~A[0] &  A[1] &  A[2] &  A[3] &  A[4] &  A[5] & ~A[6] & 
                ~A[7] & ~A[8];
assign P[ 63] =  A[0] &  A[1] &  A[2] &  A[3] &  A[4] &  A[5] & ~A[6] & 
                ~A[7] & ~A[8];
assign P[ 64] = ~A[0] & ~A[1] & ~A[2] & ~A[3] & ~A[4] & ~A[5] &  A[6] & 
                ~A[7] & ~A[8];
assign P[ 65] =  A[0] & ~A[1] & ~A[2] & ~A[3] & ~A[4] & ~A[5] &  A[6] & 
                ~A[7] & ~A[8];
assign P[ 66] = ~A[0] &  A[1] & ~A[2] & ~A[3] & ~A[4] & ~A[5] &  A[6] & 
                ~A[7] & ~A[8];
assign P[ 67] =  A[0] &  A[1] & ~A[2] & ~A[3] & ~A[4] & ~A[5] &  A[6] & 
                ~A[7] & ~A[8];
assign P[ 68] = ~A[0] & ~A[1] &  A[2] & ~A[3] & ~A[4] & ~A[5] &  A[6] & 
                ~A[7] & ~A[8];
assign P[ 69] =  A[0] & ~A[1] &  A[2] & ~A[3] & ~A[4] & ~A[5] &  A[6] & 
                ~A[7] & ~A[8];
assign P[ 70] = ~A[0] &  A[1] &  A[2] & ~A[3] & ~A[4] & ~A[5] &  A[6] & 
                ~A[7] & ~A[8];
assign P[ 71] =  A[0] &  A[1] &  A[2] & ~A[3] & ~A[4] & ~A[5] &  A[6] & 
                ~A[7] & ~A[8];
assign P[ 72] = ~A[0] & ~A[1] & ~A[2] &  A[3] & ~A[4] & ~A[5] &  A[6] & 
                ~A[7] & ~A[8];
assign P[ 73] =  A[0] & ~A[1] & ~A[2] &  A[3] & ~A[4] & ~A[5] &  A[6] & 
                ~A[7] & ~A[8];
assign P[ 74] = ~A[0] &  A[1] & ~A[2] &  A[3] & ~A[4] & ~A[5] &  A[6] & 
                ~A[7] & ~A[8];
assign P[ 75] =  A[0] &  A[1] & ~A[2] &  A[3] & ~A[4] & ~A[5] &  A[6] & 
                ~A[7] & ~A[8];
assign P[ 76] = ~A[0] & ~A[1] &  A[2] &  A[3] & ~A[4] & ~A[5] &  A[6] & 
                ~A[7] & ~A[8];
assign P[ 77] =  A[0] & ~A[1] &  A[2] &  A[3] & ~A[4] & ~A[5] &  A[6] & 
                ~A[7] & ~A[8];
assign P[ 78] = ~A[0] &  A[1] &  A[2] &  A[3] & ~A[4] & ~A[5] &  A[6] & 
                ~A[7] & ~A[8];
assign P[ 79] =  A[0] &  A[1] &  A[2] &  A[3] & ~A[4] & ~A[5] &  A[6] & 
                ~A[7] & ~A[8];
assign P[ 80] = ~A[0] & ~A[1] & ~A[2] & ~A[3] &  A[4] & ~A[5] &  A[6] & 
                ~A[7] & ~A[8];
assign P[ 81] =  A[0] & ~A[1] & ~A[2] & ~A[3] &  A[4] & ~A[5] &  A[6] & 
                ~A[7] & ~A[8];
assign P[ 82] = ~A[0] &  A[1] & ~A[2] & ~A[3] &  A[4] & ~A[5] &  A[6] & 
                ~A[7] & ~A[8];
assign P[ 83] =  A[0] &  A[1] & ~A[2] & ~A[3] &  A[4] & ~A[5] &  A[6] & 
                ~A[7] & ~A[8];
assign P[ 84] = ~A[0] & ~A[1] &  A[2] & ~A[3] &  A[4] & ~A[5] &  A[6] & 
                ~A[7] & ~A[8];
assign P[ 85] =  A[0] & ~A[1] &  A[2] & ~A[3] &  A[4] & ~A[5] &  A[6] & 
                ~A[7] & ~A[8];
assign P[ 86] = ~A[0] &  A[1] &  A[2] & ~A[3] &  A[4] & ~A[5] &  A[6] & 
                ~A[7] & ~A[8];
assign P[ 87] =  A[0] &  A[1] &  A[2] & ~A[3] &  A[4] & ~A[5] &  A[6] & 
                ~A[7] & ~A[8];
assign P[ 88] = ~A[0] & ~A[1] & ~A[2] &  A[3] &  A[4] & ~A[5] &  A[6] & 
                ~A[7] & ~A[8];
assign P[ 89] =  A[0] & ~A[1] & ~A[2] &  A[3] &  A[4] & ~A[5] &  A[6] & 
                ~A[7] & ~A[8];
assign P[ 90] = ~A[0] &  A[1] & ~A[2] &  A[3] &  A[4] & ~A[5] &  A[6] & 
                ~A[7] & ~A[8];
assign P[ 91] =  A[0] &  A[1] & ~A[2] &  A[3] &  A[4] & ~A[5] &  A[6] & 
                ~A[7] & ~A[8];
assign P[ 92] = ~A[0] & ~A[1] &  A[2] &  A[3] &  A[4] & ~A[5] &  A[6] & 
                ~A[7] & ~A[8];
assign P[ 93] =  A[0] & ~A[1] &  A[2] &  A[3] &  A[4] & ~A[5] &  A[6] & 
                ~A[7] & ~A[8];
assign P[ 94] = ~A[0] &  A[1] &  A[2] &  A[3] &  A[4] & ~A[5] &  A[6] & 
                ~A[7] & ~A[8];
assign P[ 95] =  A[0] &  A[1] &  A[2] &  A[3] &  A[4] & ~A[5] &  A[6] & 
                ~A[7] & ~A[8];
assign P[ 96] = ~A[0] & ~A[1] & ~A[2] & ~A[3] & ~A[4] &  A[5] &  A[6] & 
                ~A[7] & ~A[8];
assign P[ 97] =  A[0] & ~A[1] & ~A[2] & ~A[3] & ~A[4] &  A[5] &  A[6] & 
                ~A[7] & ~A[8];
assign P[ 98] = ~A[0] &  A[1] & ~A[2] & ~A[3] & ~A[4] &  A[5] &  A[6] & 
                ~A[7] & ~A[8];
assign P[ 99] =  A[0] &  A[1] & ~A[2] & ~A[3] & ~A[4] &  A[5] &  A[6] & 
                ~A[7] & ~A[8];
assign P[100] = ~A[0] & ~A[1] &  A[2] & ~A[3] & ~A[4] &  A[5] &  A[6] & 
                ~A[7] & ~A[8];
assign P[101] =  A[0] & ~A[1] &  A[2] & ~A[3] & ~A[4] &  A[5] &  A[6] & 
                ~A[7] & ~A[8];
assign P[102] = ~A[0] &  A[1] &  A[2] & ~A[3] & ~A[4] &  A[5] &  A[6] & 
                ~A[7] & ~A[8];
assign P[103] =  A[0] &  A[1] &  A[2] & ~A[3] & ~A[4] &  A[5] &  A[6] & 
                ~A[7] & ~A[8];
assign P[104] = ~A[0] & ~A[1] & ~A[2] &  A[3] & ~A[4] &  A[5] &  A[6] & 
                ~A[7] & ~A[8];
assign P[105] =  A[0] & ~A[1] & ~A[2] &  A[3] & ~A[4] &  A[5] &  A[6] & 
                ~A[7] & ~A[8];
assign P[106] = ~A[0] &  A[1] & ~A[2] &  A[3] & ~A[4] &  A[5] &  A[6] & 
                ~A[7] & ~A[8];
assign P[107] =  A[0] &  A[1] & ~A[2] &  A[3] & ~A[4] &  A[5] &  A[6] & 
                ~A[7] & ~A[8];
assign P[108] = ~A[0] & ~A[1] &  A[2] &  A[3] & ~A[4] &  A[5] &  A[6] & 
                ~A[7] & ~A[8];
assign P[109] =  A[0] & ~A[1] &  A[2] &  A[3] & ~A[4] &  A[5] &  A[6] & 
                ~A[7] & ~A[8];
assign P[110] = ~A[0] &  A[1] &  A[2] &  A[3] & ~A[4] &  A[5] &  A[6] & 
                ~A[7] & ~A[8];
assign P[111] =  A[0] &  A[1] &  A[2] &  A[3] & ~A[4] &  A[5] &  A[6] & 
                ~A[7] & ~A[8];
assign P[112] = ~A[0] & ~A[1] & ~A[2] & ~A[3] &  A[4] &  A[5] &  A[6] & 
                ~A[7] & ~A[8];
assign P[113] =  A[0] & ~A[1] & ~A[2] & ~A[3] &  A[4] &  A[5] &  A[6] & 
                ~A[7] & ~A[8];
assign P[114] = ~A[0] &  A[1] & ~A[2] & ~A[3] &  A[4] &  A[5] &  A[6] & 
                ~A[7] & ~A[8];
assign P[115] =  A[0] &  A[1] & ~A[2] & ~A[3] &  A[4] &  A[5] &  A[6] & 
                ~A[7] & ~A[8];
assign P[116] = ~A[0] & ~A[1] &  A[2] & ~A[3] &  A[4] &  A[5] &  A[6] & 
                ~A[7] & ~A[8];
assign P[117] =  A[0] & ~A[1] &  A[2] & ~A[3] &  A[4] &  A[5] &  A[6] & 
                ~A[7] & ~A[8];
assign P[118] = ~A[0] &  A[1] &  A[2] & ~A[3] &  A[4] &  A[5] &  A[6] & 
                ~A[7] & ~A[8];
assign P[119] =  A[0] &  A[1] &  A[2] & ~A[3] &  A[4] &  A[5] &  A[6] & 
                ~A[7] & ~A[8];
assign P[120] = ~A[0] & ~A[1] & ~A[2] &  A[3] &  A[4] &  A[5] &  A[6] & 
                ~A[7] & ~A[8];
assign P[121] =  A[0] & ~A[1] & ~A[2] &  A[3] &  A[4] &  A[5] &  A[6] & 
                ~A[7] & ~A[8];
assign P[122] = ~A[0] &  A[1] & ~A[2] &  A[3] &  A[4] &  A[5] &  A[6] & 
                ~A[7] & ~A[8];
assign P[123] =  A[0] &  A[1] & ~A[2] &  A[3] &  A[4] &  A[5] &  A[6] & 
                ~A[7] & ~A[8];
assign P[124] = ~A[0] & ~A[1] &  A[2] &  A[3] &  A[4] &  A[5] &  A[6] & 
                ~A[7] & ~A[8];
assign P[125] =  A[0] & ~A[1] &  A[2] &  A[3] &  A[4] &  A[5] &  A[6] & 
                ~A[7] & ~A[8];
assign P[126] = ~A[0] &  A[1] &  A[2] &  A[3] &  A[4] &  A[5] &  A[6] & 
                ~A[7] & ~A[8];
assign P[127] =  A[0] &  A[1] &  A[2] &  A[3] &  A[4] &  A[5] &  A[6] & 
                ~A[7] & ~A[8];
assign P[128] = ~A[0] & ~A[1] & ~A[2] & ~A[3] & ~A[4] & ~A[5] & ~A[6] & 
                 A[7] & ~A[8];
assign P[129] =  A[0] & ~A[1] & ~A[2] & ~A[3] & ~A[4] & ~A[5] & ~A[6] & 
                 A[7] & ~A[8];
assign P[130] = ~A[0] &  A[1] & ~A[2] & ~A[3] & ~A[4] & ~A[5] & ~A[6] & 
                 A[7] & ~A[8];
assign P[131] =  A[0] &  A[1] & ~A[2] & ~A[3] & ~A[4] & ~A[5] & ~A[6] & 
                 A[7] & ~A[8];
assign P[132] = ~A[0] & ~A[1] &  A[2] & ~A[3] & ~A[4] & ~A[5] & ~A[6] & 
                 A[7] & ~A[8];
assign P[133] =  A[0] & ~A[1] &  A[2] & ~A[3] & ~A[4] & ~A[5] & ~A[6] & 
                 A[7] & ~A[8];
assign P[134] = ~A[0] &  A[1] &  A[2] & ~A[3] & ~A[4] & ~A[5] & ~A[6] & 
                 A[7] & ~A[8];
assign P[135] =  A[0] &  A[1] &  A[2] & ~A[3] & ~A[4] & ~A[5] & ~A[6] & 
                 A[7] & ~A[8];
assign P[136] = ~A[0] & ~A[1] & ~A[2] &  A[3] & ~A[4] & ~A[5] & ~A[6] & 
                 A[7] & ~A[8];
assign P[137] =  A[0] & ~A[1] & ~A[2] &  A[3] & ~A[4] & ~A[5] & ~A[6] & 
                 A[7] & ~A[8];
assign P[138] = ~A[0] &  A[1] & ~A[2] &  A[3] & ~A[4] & ~A[5] & ~A[6] & 
                 A[7] & ~A[8];
assign P[139] =  A[0] &  A[1] & ~A[2] &  A[3] & ~A[4] & ~A[5] & ~A[6] & 
                 A[7] & ~A[8];
assign P[140] = ~A[0] & ~A[1] &  A[2] &  A[3] & ~A[4] & ~A[5] & ~A[6] & 
                 A[7] & ~A[8];
assign P[141] =  A[0] & ~A[1] &  A[2] &  A[3] & ~A[4] & ~A[5] & ~A[6] & 
                 A[7] & ~A[8];
assign P[142] = ~A[0] &  A[1] &  A[2] &  A[3] & ~A[4] & ~A[5] & ~A[6] & 
                 A[7] & ~A[8];
assign P[143] =  A[0] &  A[1] &  A[2] &  A[3] & ~A[4] & ~A[5] & ~A[6] & 
                 A[7] & ~A[8];
assign P[144] = ~A[0] & ~A[1] & ~A[2] & ~A[3] &  A[4] & ~A[5] & ~A[6] & 
                 A[7] & ~A[8];
assign P[145] =  A[0] & ~A[1] & ~A[2] & ~A[3] &  A[4] & ~A[5] & ~A[6] & 
                 A[7] & ~A[8];
assign P[146] = ~A[0] &  A[1] & ~A[2] & ~A[3] &  A[4] & ~A[5] & ~A[6] & 
                 A[7] & ~A[8];
assign P[147] =  A[0] &  A[1] & ~A[2] & ~A[3] &  A[4] & ~A[5] & ~A[6] & 
                 A[7] & ~A[8];
assign P[148] = ~A[0] & ~A[1] &  A[2] & ~A[3] &  A[4] & ~A[5] & ~A[6] & 
                 A[7] & ~A[8];
assign P[149] =  A[0] & ~A[1] &  A[2] & ~A[3] &  A[4] & ~A[5] & ~A[6] & 
                 A[7] & ~A[8];
assign P[150] = ~A[0] &  A[1] &  A[2] & ~A[3] &  A[4] & ~A[5] & ~A[6] & 
                 A[7] & ~A[8];
assign P[151] =  A[0] &  A[1] &  A[2] & ~A[3] &  A[4] & ~A[5] & ~A[6] & 
                 A[7] & ~A[8];
assign P[152] = ~A[0] & ~A[1] & ~A[2] &  A[3] &  A[4] & ~A[5] & ~A[6] & 
                 A[7] & ~A[8];
assign P[153] =  A[0] & ~A[1] & ~A[2] &  A[3] &  A[4] & ~A[5] & ~A[6] & 
                 A[7] & ~A[8];
assign P[154] = ~A[0] &  A[1] & ~A[2] &  A[3] &  A[4] & ~A[5] & ~A[6] & 
                 A[7] & ~A[8];
assign P[155] =  A[0] &  A[1] & ~A[2] &  A[3] &  A[4] & ~A[5] & ~A[6] & 
                 A[7] & ~A[8];
assign P[156] = ~A[0] & ~A[1] &  A[2] &  A[3] &  A[4] & ~A[5] & ~A[6] & 
                 A[7] & ~A[8];
assign P[157] =  A[0] & ~A[1] &  A[2] &  A[3] &  A[4] & ~A[5] & ~A[6] & 
                 A[7] & ~A[8];
assign P[158] = ~A[0] &  A[1] &  A[2] &  A[3] &  A[4] & ~A[5] & ~A[6] & 
                 A[7] & ~A[8];
assign P[159] =  A[0] &  A[1] &  A[2] &  A[3] &  A[4] & ~A[5] & ~A[6] & 
                 A[7] & ~A[8];
assign P[160] = ~A[0] & ~A[1] & ~A[2] & ~A[3] & ~A[4] &  A[5] & ~A[6] & 
                 A[7] & ~A[8];
assign P[161] =  A[0] & ~A[1] & ~A[2] & ~A[3] & ~A[4] &  A[5] & ~A[6] & 
                 A[7] & ~A[8];
assign P[162] = ~A[0] &  A[1] & ~A[2] & ~A[3] & ~A[4] &  A[5] & ~A[6] & 
                 A[7] & ~A[8];
assign P[163] =  A[0] &  A[1] & ~A[2] & ~A[3] & ~A[4] &  A[5] & ~A[6] & 
                 A[7] & ~A[8];
assign P[164] = ~A[0] & ~A[1] &  A[2] & ~A[3] & ~A[4] &  A[5] & ~A[6] & 
                 A[7] & ~A[8];
assign P[165] =  A[0] & ~A[1] &  A[2] & ~A[3] & ~A[4] &  A[5] & ~A[6] & 
                 A[7] & ~A[8];
assign P[166] = ~A[0] &  A[1] &  A[2] & ~A[3] & ~A[4] &  A[5] & ~A[6] & 
                 A[7] & ~A[8];
assign P[167] =  A[0] &  A[1] &  A[2] & ~A[3] & ~A[4] &  A[5] & ~A[6] & 
                 A[7] & ~A[8];
assign P[168] = ~A[0] & ~A[1] & ~A[2] &  A[3] & ~A[4] &  A[5] & ~A[6] & 
                 A[7] & ~A[8];
assign P[169] =  A[0] & ~A[1] & ~A[2] &  A[3] & ~A[4] &  A[5] & ~A[6] & 
                 A[7] & ~A[8];
assign P[170] = ~A[0] &  A[1] & ~A[2] &  A[3] & ~A[4] &  A[5] & ~A[6] & 
                 A[7] & ~A[8];
assign P[171] =  A[0] &  A[1] & ~A[2] &  A[3] & ~A[4] &  A[5] & ~A[6] & 
                 A[7] & ~A[8];
assign P[172] = ~A[0] & ~A[1] &  A[2] &  A[3] & ~A[4] &  A[5] & ~A[6] & 
                 A[7] & ~A[8];
assign P[173] =  A[0] & ~A[1] &  A[2] &  A[3] & ~A[4] &  A[5] & ~A[6] & 
                 A[7] & ~A[8];
assign P[174] = ~A[0] &  A[1] &  A[2] &  A[3] & ~A[4] &  A[5] & ~A[6] & 
                 A[7] & ~A[8];
assign P[175] =  A[0] &  A[1] &  A[2] &  A[3] & ~A[4] &  A[5] & ~A[6] & 
                 A[7] & ~A[8];
assign P[176] = ~A[0] & ~A[1] & ~A[2] & ~A[3] &  A[4] &  A[5] & ~A[6] & 
                 A[7] & ~A[8];
assign P[177] =  A[0] & ~A[1] & ~A[2] & ~A[3] &  A[4] &  A[5] & ~A[6] & 
                 A[7] & ~A[8];
assign P[178] = ~A[0] &  A[1] & ~A[2] & ~A[3] &  A[4] &  A[5] & ~A[6] & 
                 A[7] & ~A[8];
assign P[179] =  A[0] &  A[1] & ~A[2] & ~A[3] &  A[4] &  A[5] & ~A[6] & 
                 A[7] & ~A[8];
assign P[180] = ~A[0] & ~A[1] &  A[2] & ~A[3] &  A[4] &  A[5] & ~A[6] & 
                 A[7] & ~A[8];
assign P[181] =  A[0] & ~A[1] &  A[2] & ~A[3] &  A[4] &  A[5] & ~A[6] & 
                 A[7] & ~A[8];
assign P[182] = ~A[0] &  A[1] &  A[2] & ~A[3] &  A[4] &  A[5] & ~A[6] & 
                 A[7] & ~A[8];
assign P[183] =  A[0] &  A[1] &  A[2] & ~A[3] &  A[4] &  A[5] & ~A[6] & 
                 A[7] & ~A[8];
assign P[184] = ~A[0] & ~A[1] & ~A[2] &  A[3] &  A[4] &  A[5] & ~A[6] & 
                 A[7] & ~A[8];
assign P[185] =  A[0] & ~A[1] & ~A[2] &  A[3] &  A[4] &  A[5] & ~A[6] & 
                 A[7] & ~A[8];
assign P[186] = ~A[0] &  A[1] & ~A[2] &  A[3] &  A[4] &  A[5] & ~A[6] & 
                 A[7] & ~A[8];
assign P[187] =  A[0] &  A[1] & ~A[2] &  A[3] &  A[4] &  A[5] & ~A[6] & 
                 A[7] & ~A[8];
assign P[188] = ~A[0] & ~A[1] &  A[2] &  A[3] &  A[4] &  A[5] & ~A[6] & 
                 A[7] & ~A[8];
assign P[189] =  A[0] & ~A[1] &  A[2] &  A[3] &  A[4] &  A[5] & ~A[6] & 
                 A[7] & ~A[8];
assign P[190] = ~A[0] &  A[1] &  A[2] &  A[3] &  A[4] &  A[5] & ~A[6] & 
                 A[7] & ~A[8];
assign P[191] =  A[0] &  A[1] &  A[2] &  A[3] &  A[4] &  A[5] & ~A[6] & 
                 A[7] & ~A[8];
assign P[192] = ~A[0] & ~A[1] & ~A[2] & ~A[3] & ~A[4] & ~A[5] &  A[6] & 
                 A[7] & ~A[8];
assign P[193] =  A[0] & ~A[1] & ~A[2] & ~A[3] & ~A[4] & ~A[5] &  A[6] & 
                 A[7] & ~A[8];
assign P[194] = ~A[0] &  A[1] & ~A[2] & ~A[3] & ~A[4] & ~A[5] &  A[6] & 
                 A[7] & ~A[8];
assign P[195] =  A[0] &  A[1] & ~A[2] & ~A[3] & ~A[4] & ~A[5] &  A[6] & 
                 A[7] & ~A[8];
assign P[196] = ~A[0] & ~A[1] &  A[2] & ~A[3] & ~A[4] & ~A[5] &  A[6] & 
                 A[7] & ~A[8];
assign P[197] =  A[0] & ~A[1] &  A[2] & ~A[3] & ~A[4] & ~A[5] &  A[6] & 
                 A[7] & ~A[8];
assign P[198] = ~A[0] &  A[1] &  A[2] & ~A[3] & ~A[4] & ~A[5] &  A[6] & 
                 A[7] & ~A[8];
assign P[199] =  A[0] &  A[1] &  A[2] & ~A[3] & ~A[4] & ~A[5] &  A[6] & 
                 A[7] & ~A[8];
assign P[200] = ~A[0] & ~A[1] & ~A[2] &  A[3] & ~A[4] & ~A[5] &  A[6] & 
                 A[7] & ~A[8];
assign P[201] =  A[0] & ~A[1] & ~A[2] &  A[3] & ~A[4] & ~A[5] &  A[6] & 
                 A[7] & ~A[8];
assign P[202] = ~A[0] &  A[1] & ~A[2] &  A[3] & ~A[4] & ~A[5] &  A[6] & 
                 A[7] & ~A[8];
assign P[203] =  A[0] &  A[1] & ~A[2] &  A[3] & ~A[4] & ~A[5] &  A[6] & 
                 A[7] & ~A[8];
assign P[204] = ~A[0] & ~A[1] &  A[2] &  A[3] & ~A[4] & ~A[5] &  A[6] & 
                 A[7] & ~A[8];
assign P[205] =  A[0] & ~A[1] &  A[2] &  A[3] & ~A[4] & ~A[5] &  A[6] & 
                 A[7] & ~A[8];
assign P[206] = ~A[0] &  A[1] &  A[2] &  A[3] & ~A[4] & ~A[5] &  A[6] & 
                 A[7] & ~A[8];
assign P[207] =  A[0] &  A[1] &  A[2] &  A[3] & ~A[4] & ~A[5] &  A[6] & 
                 A[7] & ~A[8];
assign P[208] = ~A[0] & ~A[1] & ~A[2] & ~A[3] &  A[4] & ~A[5] &  A[6] & 
                 A[7] & ~A[8];
assign P[209] =  A[0] & ~A[1] & ~A[2] & ~A[3] &  A[4] & ~A[5] &  A[6] & 
                 A[7] & ~A[8];
assign P[210] = ~A[0] &  A[1] & ~A[2] & ~A[3] &  A[4] & ~A[5] &  A[6] & 
                 A[7] & ~A[8];
assign P[211] =  A[0] &  A[1] & ~A[2] & ~A[3] &  A[4] & ~A[5] &  A[6] & 
                 A[7] & ~A[8];
assign P[212] = ~A[0] & ~A[1] &  A[2] & ~A[3] &  A[4] & ~A[5] &  A[6] & 
                 A[7] & ~A[8];
assign P[213] =  A[0] & ~A[1] &  A[2] & ~A[3] &  A[4] & ~A[5] &  A[6] & 
                 A[7] & ~A[8];
assign P[214] = ~A[0] &  A[1] &  A[2] & ~A[3] &  A[4] & ~A[5] &  A[6] & 
                 A[7] & ~A[8];
assign P[215] =  A[0] &  A[1] &  A[2] & ~A[3] &  A[4] & ~A[5] &  A[6] & 
                 A[7] & ~A[8];
assign P[216] = ~A[0] & ~A[1] & ~A[2] &  A[3] &  A[4] & ~A[5] &  A[6] & 
                 A[7] & ~A[8];
assign P[217] =  A[0] & ~A[1] & ~A[2] &  A[3] &  A[4] & ~A[5] &  A[6] & 
                 A[7] & ~A[8];
assign P[218] = ~A[0] &  A[1] & ~A[2] &  A[3] &  A[4] & ~A[5] &  A[6] & 
                 A[7] & ~A[8];
assign P[219] =  A[0] &  A[1] & ~A[2] &  A[3] &  A[4] & ~A[5] &  A[6] & 
                 A[7] & ~A[8];
assign P[220] = ~A[0] & ~A[1] &  A[2] &  A[3] &  A[4] & ~A[5] &  A[6] & 
                 A[7] & ~A[8];
assign P[221] =  A[0] & ~A[1] &  A[2] &  A[3] &  A[4] & ~A[5] &  A[6] & 
                 A[7] & ~A[8];
assign P[222] = ~A[0] &  A[1] &  A[2] &  A[3] &  A[4] & ~A[5] &  A[6] & 
                 A[7] & ~A[8];
assign P[223] =  A[0] &  A[1] &  A[2] &  A[3] &  A[4] & ~A[5] &  A[6] & 
                 A[7] & ~A[8];
assign P[224] = ~A[0] & ~A[1] & ~A[2] & ~A[3] & ~A[4] &  A[5] &  A[6] & 
                 A[7] & ~A[8];
assign P[225] =  A[0] & ~A[1] & ~A[2] & ~A[3] & ~A[4] &  A[5] &  A[6] & 
                 A[7] & ~A[8];
assign P[226] = ~A[0] &  A[1] & ~A[2] & ~A[3] & ~A[4] &  A[5] &  A[6] & 
                 A[7] & ~A[8];
assign P[227] =  A[0] &  A[1] & ~A[2] & ~A[3] & ~A[4] &  A[5] &  A[6] & 
                 A[7] & ~A[8];
assign P[228] = ~A[0] & ~A[1] &  A[2] & ~A[3] & ~A[4] &  A[5] &  A[6] & 
                 A[7] & ~A[8];
assign P[229] =  A[0] & ~A[1] &  A[2] & ~A[3] & ~A[4] &  A[5] &  A[6] & 
                 A[7] & ~A[8];
assign P[230] = ~A[0] &  A[1] &  A[2] & ~A[3] & ~A[4] &  A[5] &  A[6] & 
                 A[7] & ~A[8];
assign P[231] =  A[0] &  A[1] &  A[2] & ~A[3] & ~A[4] &  A[5] &  A[6] & 
                 A[7] & ~A[8];
assign P[232] = ~A[0] & ~A[1] & ~A[2] &  A[3] & ~A[4] &  A[5] &  A[6] & 
                 A[7] & ~A[8];
assign P[233] =  A[0] & ~A[1] & ~A[2] &  A[3] & ~A[4] &  A[5] &  A[6] & 
                 A[7] & ~A[8];
assign P[234] = ~A[0] &  A[1] & ~A[2] &  A[3] & ~A[4] &  A[5] &  A[6] & 
                 A[7] & ~A[8];
assign P[235] =  A[0] &  A[1] & ~A[2] &  A[3] & ~A[4] &  A[5] &  A[6] & 
                 A[7] & ~A[8];
assign P[236] = ~A[0] & ~A[1] &  A[2] &  A[3] & ~A[4] &  A[5] &  A[6] & 
                 A[7] & ~A[8];
assign P[237] =  A[0] & ~A[1] &  A[2] &  A[3] & ~A[4] &  A[5] &  A[6] & 
                 A[7] & ~A[8];
assign P[238] = ~A[0] &  A[1] &  A[2] &  A[3] & ~A[4] &  A[5] &  A[6] & 
                 A[7] & ~A[8];
assign P[239] =  A[0] &  A[1] &  A[2] &  A[3] & ~A[4] &  A[5] &  A[6] & 
                 A[7] & ~A[8];
assign P[240] = ~A[0] & ~A[1] & ~A[2] & ~A[3] &  A[4] &  A[5] &  A[6] & 
                 A[7] & ~A[8];
assign P[241] =  A[0] & ~A[1] & ~A[2] & ~A[3] &  A[4] &  A[5] &  A[6] & 
                 A[7] & ~A[8];
assign P[242] = ~A[0] &  A[1] & ~A[2] & ~A[3] &  A[4] &  A[5] &  A[6] & 
                 A[7] & ~A[8];
assign P[243] =  A[0] &  A[1] & ~A[2] & ~A[3] &  A[4] &  A[5] &  A[6] & 
                 A[7] & ~A[8];
assign P[244] = ~A[0] & ~A[1] &  A[2] & ~A[3] &  A[4] &  A[5] &  A[6] & 
                 A[7] & ~A[8];
assign P[245] =  A[0] & ~A[1] &  A[2] & ~A[3] &  A[4] &  A[5] &  A[6] & 
                 A[7] & ~A[8];
assign P[246] = ~A[0] &  A[1] &  A[2] & ~A[3] &  A[4] &  A[5] &  A[6] & 
                 A[7] & ~A[8];
assign P[247] =  A[0] &  A[1] &  A[2] & ~A[3] &  A[4] &  A[5] &  A[6] & 
                 A[7] & ~A[8];
assign P[248] = ~A[0] & ~A[1] & ~A[2] &  A[3] &  A[4] &  A[5] &  A[6] & 
                 A[7] & ~A[8];
assign P[249] =  A[0] & ~A[1] & ~A[2] &  A[3] &  A[4] &  A[5] &  A[6] & 
                 A[7] & ~A[8];
assign P[250] = ~A[0] &  A[1] & ~A[2] &  A[3] &  A[4] &  A[5] &  A[6] & 
                 A[7] & ~A[8];
assign P[251] =  A[0] &  A[1] & ~A[2] &  A[3] &  A[4] &  A[5] &  A[6] & 
                 A[7] & ~A[8];
assign P[252] = ~A[0] & ~A[1] &  A[2] &  A[3] &  A[4] &  A[5] &  A[6] & 
                 A[7] & ~A[8];
assign P[253] =  A[0] & ~A[1] &  A[2] &  A[3] &  A[4] &  A[5] &  A[6] & 
                 A[7] & ~A[8];
assign P[254] = ~A[0] &  A[1] &  A[2] &  A[3] &  A[4] &  A[5] &  A[6] & 
                 A[7] & ~A[8];
assign P[255] =  A[0] &  A[1] &  A[2] &  A[3] &  A[4] &  A[5] &  A[6] & 
                 A[7] & ~A[8];
assign P[256] = ~A[0] & ~A[1] & ~A[2] & ~A[3] & ~A[4] & ~A[5] & ~A[6] & 
                ~A[7] &  A[8];
assign P[257] =  A[0] & ~A[1] & ~A[2] & ~A[3] & ~A[4] & ~A[5] & ~A[6] & 
                ~A[7] &  A[8];
assign P[258] = ~A[0] &  A[1] & ~A[2] & ~A[3] & ~A[4] & ~A[5] & ~A[6] & 
                ~A[7] &  A[8];
assign P[259] =  A[0] &  A[1] & ~A[2] & ~A[3] & ~A[4] & ~A[5] & ~A[6] & 
                ~A[7] &  A[8];
assign P[260] = ~A[0] & ~A[1] &  A[2] & ~A[3] & ~A[4] & ~A[5] & ~A[6] & 
                ~A[7] &  A[8];
assign P[261] =  A[0] & ~A[1] &  A[2] & ~A[3] & ~A[4] & ~A[5] & ~A[6] & 
                ~A[7] &  A[8];
assign P[262] = ~A[0] &  A[1] &  A[2] & ~A[3] & ~A[4] & ~A[5] & ~A[6] & 
                ~A[7] &  A[8];
assign P[263] =  A[0] &  A[1] &  A[2] & ~A[3] & ~A[4] & ~A[5] & ~A[6] & 
                ~A[7] &  A[8];
assign P[264] = ~A[0] & ~A[1] & ~A[2] &  A[3] & ~A[4] & ~A[5] & ~A[6] & 
                ~A[7] &  A[8];
assign P[265] =  A[0] & ~A[1] & ~A[2] &  A[3] & ~A[4] & ~A[5] & ~A[6] & 
                ~A[7] &  A[8];
assign P[266] = ~A[0] &  A[1] & ~A[2] &  A[3] & ~A[4] & ~A[5] & ~A[6] & 
                ~A[7] &  A[8];
assign P[267] =  A[0] &  A[1] & ~A[2] &  A[3] & ~A[4] & ~A[5] & ~A[6] & 
                ~A[7] &  A[8];
assign P[268] = ~A[0] & ~A[1] &  A[2] &  A[3] & ~A[4] & ~A[5] & ~A[6] & 
                ~A[7] &  A[8];
assign P[269] =  A[0] & ~A[1] &  A[2] &  A[3] & ~A[4] & ~A[5] & ~A[6] & 
                ~A[7] &  A[8];
assign P[270] = ~A[0] &  A[1] &  A[2] &  A[3] & ~A[4] & ~A[5] & ~A[6] & 
                ~A[7] &  A[8];
assign P[271] =  A[0] &  A[1] &  A[2] &  A[3] & ~A[4] & ~A[5] & ~A[6] & 
                ~A[7] &  A[8];
assign P[272] = ~A[0] & ~A[1] & ~A[2] & ~A[3] &  A[4] & ~A[5] & ~A[6] & 
                ~A[7] &  A[8];
assign P[273] =  A[0] & ~A[1] & ~A[2] & ~A[3] &  A[4] & ~A[5] & ~A[6] & 
                ~A[7] &  A[8];
assign P[274] = ~A[0] &  A[1] & ~A[2] & ~A[3] &  A[4] & ~A[5] & ~A[6] & 
                ~A[7] &  A[8];
assign P[275] =  A[0] &  A[1] & ~A[2] & ~A[3] &  A[4] & ~A[5] & ~A[6] & 
                ~A[7] &  A[8];
assign P[276] = ~A[0] & ~A[1] &  A[2] & ~A[3] &  A[4] & ~A[5] & ~A[6] & 
                ~A[7] &  A[8];
assign P[277] =  A[0] & ~A[1] &  A[2] & ~A[3] &  A[4] & ~A[5] & ~A[6] & 
                ~A[7] &  A[8];
assign P[278] = ~A[0] &  A[1] &  A[2] & ~A[3] &  A[4] & ~A[5] & ~A[6] & 
                ~A[7] &  A[8];
assign P[279] =  A[0] &  A[1] &  A[2] & ~A[3] &  A[4] & ~A[5] & ~A[6] & 
                ~A[7] &  A[8];
assign P[280] = ~A[0] & ~A[1] & ~A[2] &  A[3] &  A[4] & ~A[5] & ~A[6] & 
                ~A[7] &  A[8];
assign P[281] =  A[0] & ~A[1] & ~A[2] &  A[3] &  A[4] & ~A[5] & ~A[6] & 
                ~A[7] &  A[8];
assign P[282] = ~A[0] &  A[1] & ~A[2] &  A[3] &  A[4] & ~A[5] & ~A[6] & 
                ~A[7] &  A[8];
assign P[283] =  A[0] &  A[1] & ~A[2] &  A[3] &  A[4] & ~A[5] & ~A[6] & 
                ~A[7] &  A[8];
assign P[284] = ~A[0] & ~A[1] &  A[2] &  A[3] &  A[4] & ~A[5] & ~A[6] & 
                ~A[7] &  A[8];
assign P[285] =  A[0] & ~A[1] &  A[2] &  A[3] &  A[4] & ~A[5] & ~A[6] & 
                ~A[7] &  A[8];
assign P[286] = ~A[0] &  A[1] &  A[2] &  A[3] &  A[4] & ~A[5] & ~A[6] & 
                ~A[7] &  A[8];
assign P[287] =  A[0] &  A[1] &  A[2] &  A[3] &  A[4] & ~A[5] & ~A[6] & 
                ~A[7] &  A[8];
assign P[288] = ~A[0] & ~A[1] & ~A[2] & ~A[3] & ~A[4] &  A[5] & ~A[6] & 
                ~A[7] &  A[8];
assign P[289] =  A[0] & ~A[1] & ~A[2] & ~A[3] & ~A[4] &  A[5] & ~A[6] & 
                ~A[7] &  A[8];
assign P[290] = ~A[0] &  A[1] & ~A[2] & ~A[3] & ~A[4] &  A[5] & ~A[6] & 
                ~A[7] &  A[8];
assign P[291] =  A[0] &  A[1] & ~A[2] & ~A[3] & ~A[4] &  A[5] & ~A[6] & 
                ~A[7] &  A[8];
assign P[292] = ~A[0] & ~A[1] &  A[2] & ~A[3] & ~A[4] &  A[5] & ~A[6] & 
                ~A[7] &  A[8];
assign P[293] =  A[0] & ~A[1] &  A[2] & ~A[3] & ~A[4] &  A[5] & ~A[6] & 
                ~A[7] &  A[8];
assign P[294] = ~A[0] &  A[1] &  A[2] & ~A[3] & ~A[4] &  A[5] & ~A[6] & 
                ~A[7] &  A[8];
assign P[295] =  A[0] &  A[1] &  A[2] & ~A[3] & ~A[4] &  A[5] & ~A[6] & 
                ~A[7] &  A[8];
assign P[296] = ~A[0] & ~A[1] & ~A[2] &  A[3] & ~A[4] &  A[5] & ~A[6] & 
                ~A[7] &  A[8];
assign P[297] =  A[0] & ~A[1] & ~A[2] &  A[3] & ~A[4] &  A[5] & ~A[6] & 
                ~A[7] &  A[8];
assign P[298] = ~A[0] &  A[1] & ~A[2] &  A[3] & ~A[4] &  A[5] & ~A[6] & 
                ~A[7] &  A[8];
assign P[299] =  A[0] &  A[1] & ~A[2] &  A[3] & ~A[4] &  A[5] & ~A[6] & 
                ~A[7] &  A[8];
assign P[300] = ~A[0] & ~A[1] &  A[2] &  A[3] & ~A[4] &  A[5] & ~A[6] & 
                ~A[7] &  A[8];
assign P[301] =  A[0] & ~A[1] &  A[2] &  A[3] & ~A[4] &  A[5] & ~A[6] & 
                ~A[7] &  A[8];
assign P[302] = ~A[0] &  A[1] &  A[2] &  A[3] & ~A[4] &  A[5] & ~A[6] & 
                ~A[7] &  A[8];
assign P[303] =  A[0] &  A[1] &  A[2] &  A[3] & ~A[4] &  A[5] & ~A[6] & 
                ~A[7] &  A[8];
assign P[304] = ~A[0] & ~A[1] & ~A[2] & ~A[3] &  A[4] &  A[5] & ~A[6] & 
                ~A[7] &  A[8];
assign P[305] =  A[0] & ~A[1] & ~A[2] & ~A[3] &  A[4] &  A[5] & ~A[6] & 
                ~A[7] &  A[8];
assign P[306] = ~A[0] &  A[1] & ~A[2] & ~A[3] &  A[4] &  A[5] & ~A[6] & 
                ~A[7] &  A[8];
assign P[307] =  A[0] &  A[1] & ~A[2] & ~A[3] &  A[4] &  A[5] & ~A[6] & 
                ~A[7] &  A[8];
assign P[308] = ~A[0] & ~A[1] &  A[2] & ~A[3] &  A[4] &  A[5] & ~A[6] & 
                ~A[7] &  A[8];
assign P[309] =  A[0] & ~A[1] &  A[2] & ~A[3] &  A[4] &  A[5] & ~A[6] & 
                ~A[7] &  A[8];
assign P[310] = ~A[0] &  A[1] &  A[2] & ~A[3] &  A[4] &  A[5] & ~A[6] & 
                ~A[7] &  A[8];
assign P[311] =  A[0] &  A[1] &  A[2] & ~A[3] &  A[4] &  A[5] & ~A[6] & 
                ~A[7] &  A[8];
assign P[312] = ~A[0] & ~A[1] & ~A[2] &  A[3] &  A[4] &  A[5] & ~A[6] & 
                ~A[7] &  A[8];
assign P[313] =  A[0] & ~A[1] & ~A[2] &  A[3] &  A[4] &  A[5] & ~A[6] & 
                ~A[7] &  A[8];
assign P[314] = ~A[0] &  A[1] & ~A[2] &  A[3] &  A[4] &  A[5] & ~A[6] & 
                ~A[7] &  A[8];
assign P[315] =  A[0] &  A[1] & ~A[2] &  A[3] &  A[4] &  A[5] & ~A[6] & 
                ~A[7] &  A[8];
assign P[316] = ~A[0] & ~A[1] &  A[2] &  A[3] &  A[4] &  A[5] & ~A[6] & 
                ~A[7] &  A[8];
assign P[317] =  A[0] & ~A[1] &  A[2] &  A[3] &  A[4] &  A[5] & ~A[6] & 
                ~A[7] &  A[8];
assign P[318] = ~A[0] &  A[1] &  A[2] &  A[3] &  A[4] &  A[5] & ~A[6] & 
                ~A[7] &  A[8];
assign P[319] =  A[0] &  A[1] &  A[2] &  A[3] &  A[4] &  A[5] & ~A[6] & 
                ~A[7] &  A[8];
assign P[320] = ~A[0] & ~A[1] & ~A[2] & ~A[3] & ~A[4] & ~A[5] &  A[6] & 
                ~A[7] &  A[8];
assign P[321] =  A[0] & ~A[1] & ~A[2] & ~A[3] & ~A[4] & ~A[5] &  A[6] & 
                ~A[7] &  A[8];
assign P[322] = ~A[0] &  A[1] & ~A[2] & ~A[3] & ~A[4] & ~A[5] &  A[6] & 
                ~A[7] &  A[8];
assign P[323] =  A[0] &  A[1] & ~A[2] & ~A[3] & ~A[4] & ~A[5] &  A[6] & 
                ~A[7] &  A[8];
assign P[324] = ~A[0] & ~A[1] &  A[2] & ~A[3] & ~A[4] & ~A[5] &  A[6] & 
                ~A[7] &  A[8];
assign P[325] =  A[0] & ~A[1] &  A[2] & ~A[3] & ~A[4] & ~A[5] &  A[6] & 
                ~A[7] &  A[8];
assign P[326] = ~A[0] &  A[1] &  A[2] & ~A[3] & ~A[4] & ~A[5] &  A[6] & 
                ~A[7] &  A[8];
assign P[327] =  A[0] &  A[1] &  A[2] & ~A[3] & ~A[4] & ~A[5] &  A[6] & 
                ~A[7] &  A[8];
assign P[328] = ~A[0] & ~A[1] & ~A[2] &  A[3] & ~A[4] & ~A[5] &  A[6] & 
                ~A[7] &  A[8];
assign P[329] =  A[0] & ~A[1] & ~A[2] &  A[3] & ~A[4] & ~A[5] &  A[6] & 
                ~A[7] &  A[8];
assign P[330] = ~A[0] &  A[1] & ~A[2] &  A[3] & ~A[4] & ~A[5] &  A[6] & 
                ~A[7] &  A[8];
assign P[331] =  A[0] &  A[1] & ~A[2] &  A[3] & ~A[4] & ~A[5] &  A[6] & 
                ~A[7] &  A[8];
assign P[332] = ~A[0] & ~A[1] &  A[2] &  A[3] & ~A[4] & ~A[5] &  A[6] & 
                ~A[7] &  A[8];
assign P[333] =  A[0] & ~A[1] &  A[2] &  A[3] & ~A[4] & ~A[5] &  A[6] & 
                ~A[7] &  A[8];
assign P[334] = ~A[0] &  A[1] &  A[2] &  A[3] & ~A[4] & ~A[5] &  A[6] & 
                ~A[7] &  A[8];
assign P[335] =  A[0] &  A[1] &  A[2] &  A[3] & ~A[4] & ~A[5] &  A[6] & 
                ~A[7] &  A[8];
assign P[336] = ~A[0] & ~A[1] & ~A[2] & ~A[3] &  A[4] & ~A[5] &  A[6] & 
                ~A[7] &  A[8];
assign P[337] =  A[0] & ~A[1] & ~A[2] & ~A[3] &  A[4] & ~A[5] &  A[6] & 
                ~A[7] &  A[8];
assign P[338] = ~A[0] &  A[1] & ~A[2] & ~A[3] &  A[4] & ~A[5] &  A[6] & 
                ~A[7] &  A[8];
assign P[339] =  A[0] &  A[1] & ~A[2] & ~A[3] &  A[4] & ~A[5] &  A[6] & 
                ~A[7] &  A[8];
assign P[340] = ~A[0] & ~A[1] &  A[2] & ~A[3] &  A[4] & ~A[5] &  A[6] & 
                ~A[7] &  A[8];
assign P[341] =  A[0] & ~A[1] &  A[2] & ~A[3] &  A[4] & ~A[5] &  A[6] & 
                ~A[7] &  A[8];
assign P[342] = ~A[0] &  A[1] &  A[2] & ~A[3] &  A[4] & ~A[5] &  A[6] & 
                ~A[7] &  A[8];
assign P[343] =  A[0] &  A[1] &  A[2] & ~A[3] &  A[4] & ~A[5] &  A[6] & 
                ~A[7] &  A[8];
assign P[344] = ~A[0] & ~A[1] & ~A[2] &  A[3] &  A[4] & ~A[5] &  A[6] & 
                ~A[7] &  A[8];
assign P[345] =  A[0] & ~A[1] & ~A[2] &  A[3] &  A[4] & ~A[5] &  A[6] & 
                ~A[7] &  A[8];
assign P[346] = ~A[0] &  A[1] & ~A[2] &  A[3] &  A[4] & ~A[5] &  A[6] & 
                ~A[7] &  A[8];
assign P[347] =  A[0] &  A[1] & ~A[2] &  A[3] &  A[4] & ~A[5] &  A[6] & 
                ~A[7] &  A[8];
assign P[348] = ~A[0] & ~A[1] &  A[2] &  A[3] &  A[4] & ~A[5] &  A[6] & 
                ~A[7] &  A[8];
assign P[349] =  A[0] & ~A[1] &  A[2] &  A[3] &  A[4] & ~A[5] &  A[6] & 
                ~A[7] &  A[8];
assign P[350] = ~A[0] &  A[1] &  A[2] &  A[3] &  A[4] & ~A[5] &  A[6] & 
                ~A[7] &  A[8];
assign P[351] =  A[0] &  A[1] &  A[2] &  A[3] &  A[4] & ~A[5] &  A[6] & 
                ~A[7] &  A[8];
assign P[352] = ~A[0] & ~A[1] & ~A[2] & ~A[3] & ~A[4] &  A[5] &  A[6] & 
                ~A[7] &  A[8];
assign P[353] =  A[0] & ~A[1] & ~A[2] & ~A[3] & ~A[4] &  A[5] &  A[6] & 
                ~A[7] &  A[8];
assign P[354] = ~A[0] &  A[1] & ~A[2] & ~A[3] & ~A[4] &  A[5] &  A[6] & 
                ~A[7] &  A[8];
assign P[355] =  A[0] &  A[1] & ~A[2] & ~A[3] & ~A[4] &  A[5] &  A[6] & 
                ~A[7] &  A[8];
assign P[356] = ~A[0] & ~A[1] &  A[2] & ~A[3] & ~A[4] &  A[5] &  A[6] & 
                ~A[7] &  A[8];
assign P[357] =  A[0] & ~A[1] &  A[2] & ~A[3] & ~A[4] &  A[5] &  A[6] & 
                ~A[7] &  A[8];
assign P[358] = ~A[0] &  A[1] &  A[2] & ~A[3] & ~A[4] &  A[5] &  A[6] & 
                ~A[7] &  A[8];
assign P[359] =  A[0] &  A[1] &  A[2] & ~A[3] & ~A[4] &  A[5] &  A[6] & 
                ~A[7] &  A[8];
assign P[360] = ~A[0] & ~A[1] & ~A[2] &  A[3] & ~A[4] &  A[5] &  A[6] & 
                ~A[7] &  A[8];
assign P[361] =  A[0] & ~A[1] & ~A[2] &  A[3] & ~A[4] &  A[5] &  A[6] & 
                ~A[7] &  A[8];
assign P[362] = ~A[0] &  A[1] & ~A[2] &  A[3] & ~A[4] &  A[5] &  A[6] & 
                ~A[7] &  A[8];
assign P[363] =  A[0] &  A[1] & ~A[2] &  A[3] & ~A[4] &  A[5] &  A[6] & 
                ~A[7] &  A[8];
assign P[364] = ~A[0] & ~A[1] &  A[2] &  A[3] & ~A[4] &  A[5] &  A[6] & 
                ~A[7] &  A[8];
assign P[365] =  A[0] & ~A[1] &  A[2] &  A[3] & ~A[4] &  A[5] &  A[6] & 
                ~A[7] &  A[8];
assign P[366] = ~A[0] &  A[1] &  A[2] &  A[3] & ~A[4] &  A[5] &  A[6] & 
                ~A[7] &  A[8];
assign P[367] =  A[0] &  A[1] &  A[2] &  A[3] & ~A[4] &  A[5] &  A[6] & 
                ~A[7] &  A[8];
assign P[368] = ~A[0] & ~A[1] & ~A[2] & ~A[3] &  A[4] &  A[5] &  A[6] & 
                ~A[7] &  A[8];
assign P[369] =  A[0] & ~A[1] & ~A[2] & ~A[3] &  A[4] &  A[5] &  A[6] & 
                ~A[7] &  A[8];
assign P[370] = ~A[0] &  A[1] & ~A[2] & ~A[3] &  A[4] &  A[5] &  A[6] & 
                ~A[7] &  A[8];
assign P[371] =  A[0] &  A[1] & ~A[2] & ~A[3] &  A[4] &  A[5] &  A[6] & 
                ~A[7] &  A[8];
assign P[372] = ~A[0] & ~A[1] &  A[2] & ~A[3] &  A[4] &  A[5] &  A[6] & 
                ~A[7] &  A[8];
assign P[373] =  A[0] & ~A[1] &  A[2] & ~A[3] &  A[4] &  A[5] &  A[6] & 
                ~A[7] &  A[8];
assign P[374] = ~A[0] &  A[1] &  A[2] & ~A[3] &  A[4] &  A[5] &  A[6] & 
                ~A[7] &  A[8];
assign P[375] =  A[0] &  A[1] &  A[2] & ~A[3] &  A[4] &  A[5] &  A[6] & 
                ~A[7] &  A[8];
assign P[376] = ~A[0] & ~A[1] & ~A[2] &  A[3] &  A[4] &  A[5] &  A[6] & 
                ~A[7] &  A[8];
assign P[377] =  A[0] & ~A[1] & ~A[2] &  A[3] &  A[4] &  A[5] &  A[6] & 
                ~A[7] &  A[8];
assign P[378] = ~A[0] &  A[1] & ~A[2] &  A[3] &  A[4] &  A[5] &  A[6] & 
                ~A[7] &  A[8];
assign P[379] =  A[0] &  A[1] & ~A[2] &  A[3] &  A[4] &  A[5] &  A[6] & 
                ~A[7] &  A[8];
assign P[380] = ~A[0] & ~A[1] &  A[2] &  A[3] &  A[4] &  A[5] &  A[6] & 
                ~A[7] &  A[8];
assign P[381] =  A[0] & ~A[1] &  A[2] &  A[3] &  A[4] &  A[5] &  A[6] & 
                ~A[7] &  A[8];
assign P[382] = ~A[0] &  A[1] &  A[2] &  A[3] &  A[4] &  A[5] &  A[6] & 
                ~A[7] &  A[8];
assign P[383] =  A[0] &  A[1] &  A[2] &  A[3] &  A[4] &  A[5] &  A[6] & 
                ~A[7] &  A[8];
assign P[384] = ~A[0] & ~A[1] & ~A[2] & ~A[3] & ~A[4] & ~A[5] & ~A[6] & 
                 A[7] &  A[8];
assign P[385] =  A[0] & ~A[1] & ~A[2] & ~A[3] & ~A[4] & ~A[5] & ~A[6] & 
                 A[7] &  A[8];
assign P[386] = ~A[0] &  A[1] & ~A[2] & ~A[3] & ~A[4] & ~A[5] & ~A[6] & 
                 A[7] &  A[8];
assign P[387] =  A[0] &  A[1] & ~A[2] & ~A[3] & ~A[4] & ~A[5] & ~A[6] & 
                 A[7] &  A[8];
assign P[388] = ~A[0] & ~A[1] &  A[2] & ~A[3] & ~A[4] & ~A[5] & ~A[6] & 
                 A[7] &  A[8];
assign P[389] =  A[0] & ~A[1] &  A[2] & ~A[3] & ~A[4] & ~A[5] & ~A[6] & 
                 A[7] &  A[8];
assign P[390] = ~A[0] &  A[1] &  A[2] & ~A[3] & ~A[4] & ~A[5] & ~A[6] & 
                 A[7] &  A[8];
assign P[391] =  A[0] &  A[1] &  A[2] & ~A[3] & ~A[4] & ~A[5] & ~A[6] & 
                 A[7] &  A[8];
assign P[392] = ~A[0] & ~A[1] & ~A[2] &  A[3] & ~A[4] & ~A[5] & ~A[6] & 
                 A[7] &  A[8];
assign P[393] =  A[0] & ~A[1] & ~A[2] &  A[3] & ~A[4] & ~A[5] & ~A[6] & 
                 A[7] &  A[8];
assign P[394] = ~A[0] &  A[1] & ~A[2] &  A[3] & ~A[4] & ~A[5] & ~A[6] & 
                 A[7] &  A[8];
assign P[395] =  A[0] &  A[1] & ~A[2] &  A[3] & ~A[4] & ~A[5] & ~A[6] & 
                 A[7] &  A[8];
assign P[396] = ~A[0] & ~A[1] &  A[2] &  A[3] & ~A[4] & ~A[5] & ~A[6] & 
                 A[7] &  A[8];
assign P[397] =  A[0] & ~A[1] &  A[2] &  A[3] & ~A[4] & ~A[5] & ~A[6] & 
                 A[7] &  A[8];
assign P[398] = ~A[0] &  A[1] &  A[2] &  A[3] & ~A[4] & ~A[5] & ~A[6] & 
                 A[7] &  A[8];
assign P[399] =  A[0] &  A[1] &  A[2] &  A[3] & ~A[4] & ~A[5] & ~A[6] & 
                 A[7] &  A[8];
assign P[400] = ~A[0] & ~A[1] & ~A[2] & ~A[3] &  A[4] & ~A[5] & ~A[6] & 
                 A[7] &  A[8];
assign P[401] =  A[0] & ~A[1] & ~A[2] & ~A[3] &  A[4] & ~A[5] & ~A[6] & 
                 A[7] &  A[8];
assign P[402] = ~A[0] &  A[1] & ~A[2] & ~A[3] &  A[4] & ~A[5] & ~A[6] & 
                 A[7] &  A[8];
assign P[403] =  A[0] &  A[1] & ~A[2] & ~A[3] &  A[4] & ~A[5] & ~A[6] & 
                 A[7] &  A[8];
assign P[404] = ~A[0] & ~A[1] &  A[2] & ~A[3] &  A[4] & ~A[5] & ~A[6] & 
                 A[7] &  A[8];
assign P[405] =  A[0] & ~A[1] &  A[2] & ~A[3] &  A[4] & ~A[5] & ~A[6] & 
                 A[7] &  A[8];
assign P[406] = ~A[0] &  A[1] &  A[2] & ~A[3] &  A[4] & ~A[5] & ~A[6] & 
                 A[7] &  A[8];
assign P[407] =  A[0] &  A[1] &  A[2] & ~A[3] &  A[4] & ~A[5] & ~A[6] & 
                 A[7] &  A[8];
assign P[408] = ~A[0] & ~A[1] & ~A[2] &  A[3] &  A[4] & ~A[5] & ~A[6] & 
                 A[7] &  A[8];
assign P[409] =  A[0] & ~A[1] & ~A[2] &  A[3] &  A[4] & ~A[5] & ~A[6] & 
                 A[7] &  A[8];
assign P[410] = ~A[0] &  A[1] & ~A[2] &  A[3] &  A[4] & ~A[5] & ~A[6] & 
                 A[7] &  A[8];
assign P[411] =  A[0] &  A[1] & ~A[2] &  A[3] &  A[4] & ~A[5] & ~A[6] & 
                 A[7] &  A[8];
assign P[412] = ~A[0] & ~A[1] &  A[2] &  A[3] &  A[4] & ~A[5] & ~A[6] & 
                 A[7] &  A[8];
assign P[413] =  A[0] & ~A[1] &  A[2] &  A[3] &  A[4] & ~A[5] & ~A[6] & 
                 A[7] &  A[8];
assign P[414] = ~A[0] &  A[1] &  A[2] &  A[3] &  A[4] & ~A[5] & ~A[6] & 
                 A[7] &  A[8];
assign P[415] =  A[0] &  A[1] &  A[2] &  A[3] &  A[4] & ~A[5] & ~A[6] & 
                 A[7] &  A[8];
assign P[416] = ~A[0] & ~A[1] & ~A[2] & ~A[3] & ~A[4] &  A[5] & ~A[6] & 
                 A[7] &  A[8];
assign P[417] =  A[0] & ~A[1] & ~A[2] & ~A[3] & ~A[4] &  A[5] & ~A[6] & 
                 A[7] &  A[8];
assign P[418] = ~A[0] &  A[1] & ~A[2] & ~A[3] & ~A[4] &  A[5] & ~A[6] & 
                 A[7] &  A[8];
assign P[419] =  A[0] &  A[1] & ~A[2] & ~A[3] & ~A[4] &  A[5] & ~A[6] & 
                 A[7] &  A[8];
assign P[420] = ~A[0] & ~A[1] &  A[2] & ~A[3] & ~A[4] &  A[5] & ~A[6] & 
                 A[7] &  A[8];
assign P[421] =  A[0] & ~A[1] &  A[2] & ~A[3] & ~A[4] &  A[5] & ~A[6] & 
                 A[7] &  A[8];
assign P[422] = ~A[0] &  A[1] &  A[2] & ~A[3] & ~A[4] &  A[5] & ~A[6] & 
                 A[7] &  A[8];
assign P[423] =  A[0] &  A[1] &  A[2] & ~A[3] & ~A[4] &  A[5] & ~A[6] & 
                 A[7] &  A[8];
assign P[424] = ~A[0] & ~A[1] & ~A[2] &  A[3] & ~A[4] &  A[5] & ~A[6] & 
                 A[7] &  A[8];
assign P[425] =  A[0] & ~A[1] & ~A[2] &  A[3] & ~A[4] &  A[5] & ~A[6] & 
                 A[7] &  A[8];
assign P[426] = ~A[0] &  A[1] & ~A[2] &  A[3] & ~A[4] &  A[5] & ~A[6] & 
                 A[7] &  A[8];
assign P[427] =  A[0] &  A[1] & ~A[2] &  A[3] & ~A[4] &  A[5] & ~A[6] & 
                 A[7] &  A[8];
assign P[428] = ~A[0] & ~A[1] &  A[2] &  A[3] & ~A[4] &  A[5] & ~A[6] & 
                 A[7] &  A[8];
assign P[429] =  A[0] & ~A[1] &  A[2] &  A[3] & ~A[4] &  A[5] & ~A[6] & 
                 A[7] &  A[8];
assign P[430] = ~A[0] &  A[1] &  A[2] &  A[3] & ~A[4] &  A[5] & ~A[6] & 
                 A[7] &  A[8];
assign P[431] =  A[0] &  A[1] &  A[2] &  A[3] & ~A[4] &  A[5] & ~A[6] & 
                 A[7] &  A[8];
assign P[432] = ~A[0] & ~A[1] & ~A[2] & ~A[3] &  A[4] &  A[5] & ~A[6] & 
                 A[7] &  A[8];
assign P[433] =  A[0] & ~A[1] & ~A[2] & ~A[3] &  A[4] &  A[5] & ~A[6] & 
                 A[7] &  A[8];
assign P[434] = ~A[0] &  A[1] & ~A[2] & ~A[3] &  A[4] &  A[5] & ~A[6] & 
                 A[7] &  A[8];
assign P[435] =  A[0] &  A[1] & ~A[2] & ~A[3] &  A[4] &  A[5] & ~A[6] & 
                 A[7] &  A[8];
assign P[436] = ~A[0] & ~A[1] &  A[2] & ~A[3] &  A[4] &  A[5] & ~A[6] & 
                 A[7] &  A[8];
assign P[437] =  A[0] & ~A[1] &  A[2] & ~A[3] &  A[4] &  A[5] & ~A[6] & 
                 A[7] &  A[8];
assign P[438] = ~A[0] &  A[1] &  A[2] & ~A[3] &  A[4] &  A[5] & ~A[6] & 
                 A[7] &  A[8];
assign P[439] =  A[0] &  A[1] &  A[2] & ~A[3] &  A[4] &  A[5] & ~A[6] & 
                 A[7] &  A[8];
assign P[440] = ~A[0] & ~A[1] & ~A[2] &  A[3] &  A[4] &  A[5] & ~A[6] & 
                 A[7] &  A[8];
assign P[441] =  A[0] & ~A[1] & ~A[2] &  A[3] &  A[4] &  A[5] & ~A[6] & 
                 A[7] &  A[8];
assign P[442] = ~A[0] &  A[1] & ~A[2] &  A[3] &  A[4] &  A[5] & ~A[6] & 
                 A[7] &  A[8];
assign P[443] =  A[0] &  A[1] & ~A[2] &  A[3] &  A[4] &  A[5] & ~A[6] & 
                 A[7] &  A[8];
assign P[444] = ~A[0] & ~A[1] &  A[2] &  A[3] &  A[4] &  A[5] & ~A[6] & 
                 A[7] &  A[8];
assign P[445] =  A[0] & ~A[1] &  A[2] &  A[3] &  A[4] &  A[5] & ~A[6] & 
                 A[7] &  A[8];
assign P[446] = ~A[0] &  A[1] &  A[2] &  A[3] &  A[4] &  A[5] & ~A[6] & 
                 A[7] &  A[8];
assign P[447] =  A[0] &  A[1] &  A[2] &  A[3] &  A[4] &  A[5] & ~A[6] & 
                 A[7] &  A[8];
assign P[448] = ~A[0] & ~A[1] & ~A[2] & ~A[3] & ~A[4] & ~A[5] &  A[6] & 
                 A[7] &  A[8];
assign P[449] =  A[0] & ~A[1] & ~A[2] & ~A[3] & ~A[4] & ~A[5] &  A[6] & 
                 A[7] &  A[8];
assign P[450] = ~A[0] &  A[1] & ~A[2] & ~A[3] & ~A[4] & ~A[5] &  A[6] & 
                 A[7] &  A[8];
assign P[451] =  A[0] &  A[1] & ~A[2] & ~A[3] & ~A[4] & ~A[5] &  A[6] & 
                 A[7] &  A[8];
assign P[452] = ~A[0] & ~A[1] &  A[2] & ~A[3] & ~A[4] & ~A[5] &  A[6] & 
                 A[7] &  A[8];
assign P[453] =  A[0] & ~A[1] &  A[2] & ~A[3] & ~A[4] & ~A[5] &  A[6] & 
                 A[7] &  A[8];
assign P[454] = ~A[0] &  A[1] &  A[2] & ~A[3] & ~A[4] & ~A[5] &  A[6] & 
                 A[7] &  A[8];
assign P[455] =  A[0] &  A[1] &  A[2] & ~A[3] & ~A[4] & ~A[5] &  A[6] & 
                 A[7] &  A[8];
assign P[456] = ~A[0] & ~A[1] & ~A[2] &  A[3] & ~A[4] & ~A[5] &  A[6] & 
                 A[7] &  A[8];
assign P[457] =  A[0] & ~A[1] & ~A[2] &  A[3] & ~A[4] & ~A[5] &  A[6] & 
                 A[7] &  A[8];
assign P[458] = ~A[0] &  A[1] & ~A[2] &  A[3] & ~A[4] & ~A[5] &  A[6] & 
                 A[7] &  A[8];
assign P[459] =  A[0] &  A[1] & ~A[2] &  A[3] & ~A[4] & ~A[5] &  A[6] & 
                 A[7] &  A[8];
assign P[460] = ~A[0] & ~A[1] &  A[2] &  A[3] & ~A[4] & ~A[5] &  A[6] & 
                 A[7] &  A[8];
assign P[461] =  A[0] & ~A[1] &  A[2] &  A[3] & ~A[4] & ~A[5] &  A[6] & 
                 A[7] &  A[8];
assign P[462] = ~A[0] &  A[1] &  A[2] &  A[3] & ~A[4] & ~A[5] &  A[6] & 
                 A[7] &  A[8];
assign P[463] =  A[0] &  A[1] &  A[2] &  A[3] & ~A[4] & ~A[5] &  A[6] & 
                 A[7] &  A[8];
assign P[464] = ~A[0] & ~A[1] & ~A[2] & ~A[3] &  A[4] & ~A[5] &  A[6] & 
                 A[7] &  A[8];
assign P[465] =  A[0] & ~A[1] & ~A[2] & ~A[3] &  A[4] & ~A[5] &  A[6] & 
                 A[7] &  A[8];
assign P[466] = ~A[0] &  A[1] & ~A[2] & ~A[3] &  A[4] & ~A[5] &  A[6] & 
                 A[7] &  A[8];
assign P[467] =  A[0] &  A[1] & ~A[2] & ~A[3] &  A[4] & ~A[5] &  A[6] & 
                 A[7] &  A[8];
assign P[468] = ~A[0] & ~A[1] &  A[2] & ~A[3] &  A[4] & ~A[5] &  A[6] & 
                 A[7] &  A[8];
assign P[469] =  A[0] & ~A[1] &  A[2] & ~A[3] &  A[4] & ~A[5] &  A[6] & 
                 A[7] &  A[8];
assign P[470] = ~A[0] &  A[1] &  A[2] & ~A[3] &  A[4] & ~A[5] &  A[6] & 
                 A[7] &  A[8];
assign P[471] =  A[0] &  A[1] &  A[2] & ~A[3] &  A[4] & ~A[5] &  A[6] & 
                 A[7] &  A[8];
assign P[472] = ~A[0] & ~A[1] & ~A[2] &  A[3] &  A[4] & ~A[5] &  A[6] & 
                 A[7] &  A[8];
assign P[473] =  A[0] & ~A[1] & ~A[2] &  A[3] &  A[4] & ~A[5] &  A[6] & 
                 A[7] &  A[8];
assign P[474] = ~A[0] &  A[1] & ~A[2] &  A[3] &  A[4] & ~A[5] &  A[6] & 
                 A[7] &  A[8];
assign P[475] =  A[0] &  A[1] & ~A[2] &  A[3] &  A[4] & ~A[5] &  A[6] & 
                 A[7] &  A[8];
assign P[476] = ~A[0] & ~A[1] &  A[2] &  A[3] &  A[4] & ~A[5] &  A[6] & 
                 A[7] &  A[8];
assign P[477] =  A[0] & ~A[1] &  A[2] &  A[3] &  A[4] & ~A[5] &  A[6] & 
                 A[7] &  A[8];
assign P[478] = ~A[0] &  A[1] &  A[2] &  A[3] &  A[4] & ~A[5] &  A[6] & 
                 A[7] &  A[8];
assign P[479] =  A[0] &  A[1] &  A[2] &  A[3] &  A[4] & ~A[5] &  A[6] & 
                 A[7] &  A[8];
assign P[480] = ~A[0] & ~A[1] & ~A[2] & ~A[3] & ~A[4] &  A[5] &  A[6] & 
                 A[7] &  A[8];
assign P[481] =  A[0] & ~A[1] & ~A[2] & ~A[3] & ~A[4] &  A[5] &  A[6] & 
                 A[7] &  A[8];
assign P[482] = ~A[0] &  A[1] & ~A[2] & ~A[3] & ~A[4] &  A[5] &  A[6] & 
                 A[7] &  A[8];
assign P[483] =  A[0] &  A[1] & ~A[2] & ~A[3] & ~A[4] &  A[5] &  A[6] & 
                 A[7] &  A[8];
assign P[484] = ~A[0] & ~A[1] &  A[2] & ~A[3] & ~A[4] &  A[5] &  A[6] & 
                 A[7] &  A[8];
assign P[485] =  A[0] & ~A[1] &  A[2] & ~A[3] & ~A[4] &  A[5] &  A[6] & 
                 A[7] &  A[8];
assign P[486] = ~A[0] &  A[1] &  A[2] & ~A[3] & ~A[4] &  A[5] &  A[6] & 
                 A[7] &  A[8];
assign P[487] =  A[0] &  A[1] &  A[2] & ~A[3] & ~A[4] &  A[5] &  A[6] & 
                 A[7] &  A[8];
assign P[488] = ~A[0] & ~A[1] & ~A[2] &  A[3] & ~A[4] &  A[5] &  A[6] & 
                 A[7] &  A[8];
assign P[489] =  A[0] & ~A[1] & ~A[2] &  A[3] & ~A[4] &  A[5] &  A[6] & 
                 A[7] &  A[8];
assign P[490] = ~A[0] &  A[1] & ~A[2] &  A[3] & ~A[4] &  A[5] &  A[6] & 
                 A[7] &  A[8];
assign P[491] =  A[0] &  A[1] & ~A[2] &  A[3] & ~A[4] &  A[5] &  A[6] & 
                 A[7] &  A[8];
assign P[492] = ~A[0] & ~A[1] &  A[2] &  A[3] & ~A[4] &  A[5] &  A[6] & 
                 A[7] &  A[8];
assign P[493] =  A[0] & ~A[1] &  A[2] &  A[3] & ~A[4] &  A[5] &  A[6] & 
                 A[7] &  A[8];
assign P[494] = ~A[0] &  A[1] &  A[2] &  A[3] & ~A[4] &  A[5] &  A[6] & 
                 A[7] &  A[8];
assign P[495] =  A[0] &  A[1] &  A[2] &  A[3] & ~A[4] &  A[5] &  A[6] & 
                 A[7] &  A[8];
assign P[496] = ~A[0] & ~A[1] & ~A[2] & ~A[3] &  A[4] &  A[5] &  A[6] & 
                 A[7] &  A[8];
assign P[497] =  A[0] & ~A[1] & ~A[2] & ~A[3] &  A[4] &  A[5] &  A[6] & 
                 A[7] &  A[8];
assign P[498] = ~A[0] &  A[1] & ~A[2] & ~A[3] &  A[4] &  A[5] &  A[6] & 
                 A[7] &  A[8];
assign P[499] =  A[0] &  A[1] & ~A[2] & ~A[3] &  A[4] &  A[5] &  A[6] & 
                 A[7] &  A[8];
assign P[500] = ~A[0] & ~A[1] &  A[2] & ~A[3] &  A[4] &  A[5] &  A[6] & 
                 A[7] &  A[8];
assign P[501] =  A[0] & ~A[1] &  A[2] & ~A[3] &  A[4] &  A[5] &  A[6] & 
                 A[7] &  A[8];
assign P[502] = ~A[0] &  A[1] &  A[2] & ~A[3] &  A[4] &  A[5] &  A[6] & 
                 A[7] &  A[8];
assign P[503] =  A[0] &  A[1] &  A[2] & ~A[3] &  A[4] &  A[5] &  A[6] & 
                 A[7] &  A[8];
assign P[504] = ~A[0] & ~A[1] & ~A[2] &  A[3] &  A[4] &  A[5] &  A[6] & 
                 A[7] &  A[8];
assign P[505] =  A[0] & ~A[1] & ~A[2] &  A[3] &  A[4] &  A[5] &  A[6] & 
                 A[7] &  A[8];
assign P[506] = ~A[0] &  A[1] & ~A[2] &  A[3] &  A[4] &  A[5] &  A[6] & 
                 A[7] &  A[8];
assign P[507] =  A[0] &  A[1] & ~A[2] &  A[3] &  A[4] &  A[5] &  A[6] & 
                 A[7] &  A[8];
assign P[508] = ~A[0] & ~A[1] &  A[2] &  A[3] &  A[4] &  A[5] &  A[6] & 
                 A[7] &  A[8];
assign P[509] =  A[0] & ~A[1] &  A[2] &  A[3] &  A[4] &  A[5] &  A[6] & 
                 A[7] &  A[8];
assign P[510] = ~A[0] &  A[1] &  A[2] &  A[3] &  A[4] &  A[5] &  A[6] & 
                 A[7] &  A[8];
assign P[511] =  A[0] &  A[1] &  A[2] &  A[3] &  A[4] &  A[5] &  A[6] & 
                 A[7] &  A[8];

always @(posedge Clk)
begin
    if(Rst)
        Q <= #1 0;
    else if(CE) begin
        Q[ 0] <= #1 P[183] | P[192] | P[193] | P[207] | P[439];
        Q[ 1] <= #1 P[183] | P[184] | P[185] | P[194] | P[195] | P[196] | 
                    P[197] | P[198] | P[199] | P[200] | P[201] | P[202] | 
                    P[203] | P[204] | P[205] | P[208] | P[435] | P[437] | 
                    P[439];
        Q[ 2] <= #1 P[183] | P[186] | P[188] | P[192] | P[193] | P[208];
        Q[ 3] <= #1 P[  3] | P[  5] | P[ 12] | P[ 14];
        Q[ 4] <= #1 P[  1] | P[  2] | P[  3] | P[  8] | P[  9] | P[ 10] | 
                    P[ 11] | P[ 12] | P[ 24] | P[ 39] | P[ 40] | P[ 42] | 
                    P[ 43] | P[ 45] | P[ 46] | P[ 47] | P[ 70] | P[ 71] | 
                    P[ 76] | P[ 77] | P[ 82] | P[ 83] | P[102] | P[103] | 
                    P[107] | P[108] | P[112] | P[113] | P[121] | P[129] | 
                    P[132] | P[133] | P[135] | P[139] | P[143] | P[151] | 
                    P[152] | P[154] | P[155] | P[157] | P[158] | P[165] | 
                    P[169] | P[178] | P[181] | P[182] | P[183] | P[190] | 
                    P[193] | P[200] | P[201] | P[206] | P[207] | P[208] | 
                    P[214] | P[217] | P[218] | P[220] | P[384] | P[385] | 
                    P[387] | P[388] | P[389] | P[391] | P[392] | P[393] | 
                    P[394] | P[395] | P[396] | P[397] | P[398] | P[399] | 
                    P[416] | P[417] | P[418] | P[419] | P[420] | P[421] | 
                    P[422] | P[424] | P[425] | P[426] | P[427] | P[428] | 
                    P[429] | P[432] | P[433] | P[434] | P[436] | P[439];
        Q[ 5] <= #1 P[ 47] | P[ 70] | P[ 71] | P[ 76] | P[ 77] | P[ 82] | 
                    P[ 83] | P[102] | P[103] | P[107] | P[108] | P[112] | 
                    P[113] | P[121] | P[129] | P[132] | P[133] | P[135] | 
                    P[139] | P[143] | P[157] | P[158] | P[165] | P[169] | 
                    P[178] | P[181] | P[182] | P[183] | P[190] | P[200] | 
                    P[201] | P[206] | P[208] | P[214] | P[217] | P[218] | 
                    P[220] | P[257] | P[259] | P[261] | P[263] | P[264] | 
                    P[265] | P[267] | P[269] | P[271] | P[272] | P[274] | 
                    P[276] | P[278] | P[280] | P[282] | P[284] | P[286] | 
                    P[300] | P[304] | P[305] | P[306] | P[307] | P[308] | 
                    P[309] | P[310] | P[311] | P[312] | P[313] | P[314] | 
                    P[315] | P[316] | P[317] | P[318] | P[319] | P[323] | 
                    P[324] | P[327] | P[329] | P[331] | P[337] | P[339] | 
                    P[341] | P[343] | P[345] | P[347] | P[349] | P[351] | 
                    P[353] | P[355] | P[357] | P[359] | P[365] | P[367] | 
                    P[384] | P[388] | P[421] | P[429] | P[436] | P[439];
        Q[ 6] <= #1 P[  1] | P[  4] | P[  5] | P[  9] | P[ 10] | P[ 13] | 
                    P[ 14] | P[ 16] | P[ 18] | P[ 19] | P[ 21] | P[ 22] | 
                    P[ 24] | P[ 25] | P[ 27] | P[ 28] | P[ 29] | P[ 30] | 
                    P[ 31] | P[ 32] | P[ 33] | P[ 34] | P[ 35] | P[ 36] | 
                    P[ 37] | P[ 40] | P[ 41] | P[ 43] | P[ 44] | P[ 46] | 
                    P[ 48] | P[ 49] | P[ 50] | P[ 51] | P[ 52] | P[ 53] | 
                    P[ 54] | P[ 55] | P[ 56] | P[ 57] | P[ 58] | P[ 59] | 
                    P[ 60] | P[ 61] | P[ 62] | P[ 63] | P[ 64] | P[ 65] | 
                    P[ 66] | P[ 67] | P[ 68] | P[ 69] | P[ 72] | P[ 73] | 
                    P[ 74] | P[ 75] | P[ 78] | P[ 79] | P[ 80] | P[ 81] | 
                    P[ 84] | P[ 85] | P[ 86] | P[ 87] | P[ 88] | P[ 89] | 
                    P[ 90] | P[ 91] | P[ 92] | P[ 93] | P[ 94] | P[ 95] | 
                    P[ 96] | P[ 97] | P[ 98] | P[ 99] | P[100] | P[101] | 
                    P[104] | P[105] | P[106] | P[109] | P[110] | P[111] | 
                    P[115] | P[116] | P[117] | P[118] | P[119] | P[120] | 
                    P[122] | P[123] | P[124] | P[125] | P[126] | P[127] | 
                    P[128] | P[130] | P[131] | P[134] | P[136] | P[137] | 
                    P[138] | P[140] | P[141] | P[142] | P[143] | P[149] | 
                    P[151] | P[154] | P[156] | P[157] | P[159] | P[160] | 
                    P[161] | P[162] | P[163] | P[164] | P[166] | P[167] | 
                    P[168] | P[169] | P[170] | P[171] | P[173] | P[174] | 
                    P[175] | P[177] | P[179] | P[180] | P[182] | P[184] | 
                    P[185] | P[186] | P[187] | P[191] | P[193] | P[194] | 
                    P[195] | P[196] | P[197] | P[198] | P[199] | P[202] | 
                    P[203] | P[204] | P[205] | P[210] | P[211] | P[212] | 
                    P[213] | P[215] | P[216] | P[219] | P[256] | P[257] | 
                    P[258] | P[259] | P[260] | P[261] | P[262] | P[263] | 
                    P[264] | P[265] | P[266] | P[267] | P[268] | P[269] | 
                    P[270] | P[271] | P[272] | P[273] | P[274] | P[275] | 
                    P[276] | P[277] | P[278] | P[279] | P[280] | P[281] | 
                    P[282] | P[283] | P[284] | P[285] | P[286] | P[287] | 
                    P[288] | P[289] | P[291] | P[293] | P[295] | P[297] | 
                    P[298] | P[299] | P[300] | P[301] | P[302] | P[303] | 
                    P[304] | P[305] | P[306] | P[307] | P[308] | P[309] | 
                    P[310] | P[311] | P[312] | P[313] | P[314] | P[315] | 
                    P[316] | P[317] | P[318] | P[319] | P[320] | P[321] | 
                    P[322] | P[323] | P[324] | P[325] | P[326] | P[327] | 
                    P[328] | P[329] | P[330] | P[331] | P[332] | P[333] | 
                    P[334] | P[335] | P[336] | P[337] | P[338] | P[339] | 
                    P[340] | P[341] | P[342] | P[343] | P[344] | P[345] | 
                    P[346] | P[347] | P[348] | P[349] | P[350] | P[351] | 
                    P[352] | P[353] | P[354] | P[355] | P[356] | P[357] | 
                    P[358] | P[359] | P[360] | P[361] | P[362] | P[363] | 
                    P[364] | P[365] | P[366] | P[367] | P[368] | P[369] | 
                    P[370] | P[371] | P[372] | P[373] | P[374] | P[375] | 
                    P[376] | P[377] | P[378] | P[379] | P[380] | P[381] | 
                    P[382] | P[383] | P[386] | P[390] | P[400] | P[401] | 
                    P[402] | P[403] | P[404] | P[405] | P[406] | P[407] | 
                    P[408] | P[409] | P[410] | P[411] | P[412] | P[413] | 
                    P[414] | P[415] | P[423] | P[431] | P[435] | P[436] | 
                    P[438] | P[439] | P[448] | P[449] | P[450] | P[451] | 
                    P[452] | P[453] | P[454] | P[455] | P[456] | P[457] | 
                    P[458] | P[459] | P[460] | P[461] | P[462] | P[463] | 
                    P[464] | P[465] | P[466] | P[467] | P[468] | P[469] | 
                    P[470] | P[471] | P[472] | P[473] | P[474] | P[475] | 
                    P[476] | P[477] | P[478] | P[479] | P[480] | P[481] | 
                    P[482] | P[483] | P[484] | P[485] | P[486] | P[487] | 
                    P[488] | P[489] | P[490] | P[491] | P[492] | P[493] | 
                    P[494] | P[495] | P[496] | P[497] | P[498] | P[499] | 
                    P[500] | P[501] | P[502] | P[503] | P[504] | P[505] | 
                    P[506] | P[507] | P[508] | P[509] | P[510] | P[511];
        Q[ 7] <= #1 P[  2] | P[  4] | P[ 11] | P[ 13] | P[ 20] | P[ 21] | 
                    P[ 24] | P[ 28] | P[ 30] | P[ 34] | P[ 36] | P[ 48] | 
                    P[ 50] | P[ 52] | P[ 54] | P[ 56] | P[ 58] | P[ 60] | 
                    P[ 62] | P[ 64] | P[ 66] | P[ 68] | P[ 72] | P[ 74] | 
                    P[ 78] | P[ 80] | P[ 85] | P[ 87] | P[ 90] | P[ 92] | 
                    P[ 95] | P[ 97] | P[100] | P[105] | P[110] | P[116] | 
                    P[117] | P[123] | P[125] | P[130] | P[134] | P[136] | 
                    P[138] | P[140] | P[142] | P[143] | P[152] | P[155] | 
                    P[158] | P[159] | P[161] | P[165] | P[166] | P[167] | 
                    P[170] | P[174] | P[177] | P[178] | P[179] | P[181] | 
                    P[183] | P[184] | P[186] | P[190] | P[194] | P[196] | 
                    P[198] | P[202] | P[207] | P[210] | P[215] | P[219] | 
                    P[256] | P[257] | P[258] | P[259] | P[260] | P[261] | 
                    P[262] | P[263] | P[264] | P[265] | P[266] | P[267] | 
                    P[268] | P[269] | P[270] | P[271] | P[272] | P[273] | 
                    P[274] | P[275] | P[276] | P[277] | P[278] | P[279] | 
                    P[280] | P[281] | P[282] | P[283] | P[284] | P[285] | 
                    P[286] | P[287] | P[289] | P[291] | P[293] | P[295] | 
                    P[297] | P[298] | P[299] | P[300] | P[301] | P[302] | 
                    P[303] | P[304] | P[305] | P[306] | P[307] | P[308] | 
                    P[309] | P[310] | P[311] | P[312] | P[313] | P[314] | 
                    P[315] | P[316] | P[317] | P[318] | P[319] | P[320] | 
                    P[321] | P[322] | P[323] | P[324] | P[326] | P[327] | 
                    P[328] | P[329] | P[330] | P[331] | P[332] | P[333] | 
                    P[334] | P[335] | P[336] | P[337] | P[338] | P[339] | 
                    P[340] | P[341] | P[342] | P[343] | P[344] | P[345] | 
                    P[346] | P[347] | P[348] | P[349] | P[350] | P[351] | 
                    P[352] | P[353] | P[354] | P[355] | P[356] | P[357] | 
                    P[358] | P[359] | P[360] | P[361] | P[362] | P[363] | 
                    P[364] | P[365] | P[366] | P[367] | P[368] | P[369] | 
                    P[370] | P[371] | P[372] | P[373] | P[374] | P[375] | 
                    P[376] | P[377] | P[378] | P[379] | P[380] | P[381] | 
                    P[382] | P[383] | P[386] | P[390] | P[400] | P[401] | 
                    P[402] | P[403] | P[404] | P[405] | P[406] | P[407] | 
                    P[408] | P[409] | P[410] | P[411] | P[412] | P[413] | 
                    P[414] | P[415] | P[423] | P[431] | P[435] | P[438] | 
                    P[448] | P[449] | P[450] | P[451] | P[452] | P[453] | 
                    P[454] | P[455] | P[456] | P[457] | P[458] | P[459] | 
                    P[460] | P[461] | P[462] | P[463] | P[464] | P[465] | 
                    P[466] | P[467] | P[468] | P[469] | P[470] | P[471] | 
                    P[472] | P[473] | P[474] | P[475] | P[476] | P[477] | 
                    P[478] | P[479] | P[480] | P[481] | P[482] | P[483] | 
                    P[484] | P[485] | P[486] | P[487] | P[488] | P[489] | 
                    P[490] | P[491] | P[492] | P[493] | P[494] | P[495] | 
                    P[496] | P[497] | P[498] | P[499] | P[500] | P[501] | 
                    P[502] | P[503] | P[504] | P[505] | P[506] | P[507] | 
                    P[508] | P[509] | P[510] | P[511];
        Q[ 8] <= #1 P[  3] | P[  6] | P[  8] | P[ 12] | P[ 15] | P[ 17] | 
                    P[ 23] | P[ 26] | P[ 38] | P[ 39] | P[ 42] | P[ 45] | 
                    P[114] | P[144] | P[153] | P[188] | P[189] | P[192] | 
                    P[209] | P[290] | P[292] | P[294] | P[296] | P[385] | 
                    P[387] | P[389] | P[391] | P[392] | P[393] | P[394] | 
                    P[395] | P[396] | P[397] | P[398] | P[399] | P[416] | 
                    P[417] | P[418] | P[419] | P[420] | P[422] | P[424] | 
                    P[425] | P[426] | P[427] | P[428] | P[430] | P[432] | 
                    P[433] | P[434] | P[437] | P[440] | P[441] | P[442] | 
                    P[443] | P[444] | P[445] | P[446] | P[447];
        Q[ 9] <= #1 P[  1] | P[  2] | P[  3] | P[  9] | P[ 10] | P[ 11] | 
                    P[ 12] | P[ 19] | P[ 20] | P[ 40] | P[ 43] | P[ 46] | 
                    P[ 47] | P[ 70] | P[ 71] | P[ 76] | P[ 77] | P[ 82] | 
                    P[ 83] | P[102] | P[103] | P[107] | P[108] | P[112] | 
                    P[113] | P[115] | P[121] | P[129] | P[132] | P[133] | 
                    P[135] | P[139] | P[151] | P[152] | P[154] | P[155] | 
                    P[157] | P[158] | P[165] | P[169] | P[178] | P[181] | 
                    P[182] | P[183] | P[190] | P[193] | P[200] | P[201] | 
                    P[206] | P[208] | P[214] | P[217] | P[218] | P[220] | 
                    P[384] | P[388] | P[421] | P[429] | P[436] | P[439];
        Q[10] <= #1 P[  4] | P[  5] | P[  6] | P[  8] | P[ 13] | P[ 14] | 
                    P[ 15] | P[ 16] | P[ 17] | P[ 18] | P[ 21] | P[ 22] | 
                    P[ 23] | P[ 24] | P[ 25] | P[ 26] | P[ 27] | P[ 28] | 
                    P[ 29] | P[ 30] | P[ 31] | P[ 32] | P[ 33] | P[ 34] | 
                    P[ 35] | P[ 36] | P[ 37] | P[ 38] | P[ 39] | P[ 41] | 
                    P[ 42] | P[ 44] | P[ 45] | P[ 48] | P[ 49] | P[ 50] | 
                    P[ 51] | P[ 52] | P[ 53] | P[ 54] | P[ 55] | P[ 56] | 
                    P[ 57] | P[ 58] | P[ 59] | P[ 60] | P[ 61] | P[ 62] | 
                    P[ 63] | P[ 64] | P[ 65] | P[ 66] | P[ 67] | P[ 68] | 
                    P[ 69] | P[ 72] | P[ 73] | P[ 74] | P[ 75] | P[ 78] | 
                    P[ 79] | P[ 80] | P[ 81] | P[ 84] | P[ 85] | P[ 86] | 
                    P[ 87] | P[ 88] | P[ 89] | P[ 90] | P[ 91] | P[ 92] | 
                    P[ 93] | P[ 94] | P[ 95] | P[ 96] | P[ 97] | P[ 98] | 
                    P[ 99] | P[100] | P[101] | P[104] | P[105] | P[106] | 
                    P[109] | P[110] | P[111] | P[114] | P[116] | P[117] | 
                    P[118] | P[119] | P[120] | P[122] | P[123] | P[124] | 
                    P[125] | P[126] | P[127] | P[128] | P[130] | P[131] | 
                    P[134] | P[136] | P[137] | P[138] | P[140] | P[141] | 
                    P[142] | P[143] | P[144] | P[149] | P[153] | P[156] | 
                    P[159] | P[160] | P[161] | P[162] | P[163] | P[164] | 
                    P[166] | P[167] | P[168] | P[170] | P[171] | P[173] | 
                    P[174] | P[175] | P[177] | P[179] | P[180] | P[184] | 
                    P[185] | P[186] | P[187] | P[188] | P[189] | P[191] | 
                    P[192] | P[194] | P[195] | P[196] | P[197] | P[198] | 
                    P[199] | P[202] | P[203] | P[204] | P[205] | P[207] | 
                    P[209] | P[210] | P[211] | P[212] | P[213] | P[215] | 
                    P[216] | P[219] | P[256] | P[257] | P[258] | P[259] | 
                    P[260] | P[261] | P[262] | P[263] | P[264] | P[265] | 
                    P[266] | P[267] | P[268] | P[269] | P[270] | P[271] | 
                    P[272] | P[273] | P[274] | P[275] | P[276] | P[277] | 
                    P[278] | P[279] | P[280] | P[281] | P[282] | P[283] | 
                    P[284] | P[285] | P[286] | P[287] | P[288] | P[289] | 
                    P[290] | P[291] | P[292] | P[293] | P[294] | P[295] | 
                    P[296] | P[297] | P[298] | P[299] | P[300] | P[301] | 
                    P[302] | P[303] | P[304] | P[305] | P[306] | P[307] | 
                    P[308] | P[309] | P[310] | P[311] | P[312] | P[313] | 
                    P[314] | P[315] | P[316] | P[317] | P[318] | P[319] | 
                    P[320] | P[321] | P[322] | P[323] | P[324] | P[325] | 
                    P[326] | P[327] | P[328] | P[329] | P[330] | P[331] | 
                    P[332] | P[333] | P[334] | P[335] | P[336] | P[337] | 
                    P[338] | P[339] | P[340] | P[341] | P[342] | P[343] | 
                    P[344] | P[345] | P[346] | P[347] | P[348] | P[349] | 
                    P[350] | P[351] | P[352] | P[353] | P[354] | P[355] | 
                    P[356] | P[357] | P[358] | P[359] | P[360] | P[361] | 
                    P[362] | P[363] | P[364] | P[365] | P[366] | P[367] | 
                    P[368] | P[369] | P[370] | P[371] | P[372] | P[373] | 
                    P[374] | P[375] | P[376] | P[377] | P[378] | P[379] | 
                    P[380] | P[381] | P[382] | P[383] | P[385] | P[386] | 
                    P[387] | P[389] | P[390] | P[391] | P[392] | P[393] | 
                    P[394] | P[395] | P[396] | P[397] | P[398] | P[399] | 
                    P[400] | P[401] | P[402] | P[403] | P[404] | P[405] | 
                    P[406] | P[407] | P[408] | P[409] | P[410] | P[411] | 
                    P[412] | P[413] | P[414] | P[415] | P[416] | P[417] | 
                    P[418] | P[419] | P[420] | P[422] | P[423] | P[424] | 
                    P[425] | P[426] | P[427] | P[428] | P[430] | P[431] | 
                    P[432] | P[433] | P[434] | P[435] | P[437] | P[438] | 
                    P[440] | P[441] | P[442] | P[443] | P[444] | P[445] | 
                    P[446] | P[447] | P[448] | P[449] | P[450] | P[451] | 
                    P[452] | P[453] | P[454] | P[455] | P[456] | P[457] | 
                    P[458] | P[459] | P[460] | P[461] | P[462] | P[463] | 
                    P[464] | P[465] | P[466] | P[467] | P[468] | P[469] | 
                    P[470] | P[471] | P[472] | P[473] | P[474] | P[475] | 
                    P[476] | P[477] | P[478] | P[479] | P[480] | P[481] | 
                    P[482] | P[483] | P[484] | P[485] | P[486] | P[487] | 
                    P[488] | P[489] | P[490] | P[491] | P[492] | P[493] | 
                    P[494] | P[495] | P[496] | P[497] | P[498] | P[499] | 
                    P[500] | P[501] | P[502] | P[503] | P[504] | P[505] | 
                    P[506] | P[507] | P[508] | P[509] | P[510] | P[511];
        Q[11] <= #1 P[  5] | P[  8] | P[ 14] | P[ 16] | P[ 17] | P[ 18] | 
                    P[ 22] | P[ 24] | P[ 25] | P[ 26] | P[ 27] | P[ 29] | 
                    P[ 31] | P[ 32] | P[ 33] | P[ 35] | P[ 37] | P[ 39] | 
                    P[ 41] | P[ 42] | P[ 44] | P[ 45] | P[ 49] | P[ 51] | 
                    P[ 53] | P[ 55] | P[ 57] | P[ 59] | P[ 61] | P[ 63] | 
                    P[ 65] | P[ 67] | P[ 69] | P[ 71] | P[ 73] | P[ 75] | 
                    P[ 77] | P[ 79] | P[ 81] | P[ 83] | P[ 84] | P[ 86] | 
                    P[ 88] | P[ 89] | P[ 91] | P[ 93] | P[ 94] | P[ 96] | 
                    P[ 98] | P[ 99] | P[101] | P[103] | P[104] | P[106] | 
                    P[108] | P[109] | P[111] | P[113] | P[114] | P[118] | 
                    P[119] | P[120] | P[122] | P[124] | P[126] | P[127] | 
                    P[128] | P[131] | P[133] | P[137] | P[141] | P[143] | 
                    P[144] | P[149] | P[150] | P[153] | P[156] | P[160] | 
                    P[162] | P[163] | P[164] | P[168] | P[171] | P[173] | 
                    P[175] | P[177] | P[179] | P[180] | P[182] | P[187] | 
                    P[191] | P[192] | P[203] | P[204] | P[205] | P[209] | 
                    P[211] | P[212] | P[213] | P[216] | P[218] | P[256] | 
                    P[257] | P[258] | P[259] | P[260] | P[261] | P[262] | 
                    P[263] | P[264] | P[265] | P[266] | P[267] | P[268] | 
                    P[269] | P[270] | P[271] | P[272] | P[273] | P[274] | 
                    P[275] | P[276] | P[277] | P[278] | P[279] | P[280] | 
                    P[281] | P[282] | P[283] | P[284] | P[285] | P[286] | 
                    P[287] | P[288] | P[289] | P[290] | P[291] | P[292] | 
                    P[293] | P[294] | P[295] | P[296] | P[297] | P[298] | 
                    P[299] | P[300] | P[301] | P[302] | P[303] | P[304] | 
                    P[305] | P[306] | P[307] | P[308] | P[309] | P[310] | 
                    P[311] | P[312] | P[313] | P[314] | P[315] | P[316] | 
                    P[317] | P[318] | P[319] | P[320] | P[321] | P[322] | 
                    P[323] | P[324] | P[325] | P[326] | P[327] | P[328] | 
                    P[329] | P[330] | P[331] | P[332] | P[333] | P[334] | 
                    P[335] | P[336] | P[337] | P[338] | P[339] | P[340] | 
                    P[341] | P[342] | P[343] | P[344] | P[345] | P[346] | 
                    P[347] | P[348] | P[349] | P[350] | P[351] | P[352] | 
                    P[353] | P[354] | P[355] | P[356] | P[357] | P[358] | 
                    P[359] | P[360] | P[361] | P[362] | P[363] | P[364] | 
                    P[365] | P[366] | P[367] | P[368] | P[369] | P[370] | 
                    P[371] | P[372] | P[373] | P[374] | P[375] | P[376] | 
                    P[377] | P[378] | P[379] | P[380] | P[381] | P[382] | 
                    P[383] | P[385] | P[386] | P[387] | P[389] | P[390] | 
                    P[391] | P[392] | P[393] | P[394] | P[395] | P[396] | 
                    P[397] | P[398] | P[399] | P[400] | P[401] | P[402] | 
                    P[403] | P[404] | P[405] | P[406] | P[407] | P[408] | 
                    P[409] | P[410] | P[411] | P[412] | P[413] | P[414] | 
                    P[415] | P[416] | P[417] | P[418] | P[419] | P[420] | 
                    P[422] | P[423] | P[424] | P[425] | P[426] | P[427] | 
                    P[428] | P[430] | P[431] | P[432] | P[433] | P[434] | 
                    P[437] | P[438] | P[440] | P[441] | P[442] | P[443] | 
                    P[444] | P[445] | P[446] | P[447] | P[448] | P[449] | 
                    P[450] | P[451] | P[452] | P[453] | P[454] | P[455] | 
                    P[456] | P[457] | P[458] | P[459] | P[460] | P[461] | 
                    P[462] | P[463] | P[464] | P[465] | P[466] | P[467] | 
                    P[468] | P[469] | P[470] | P[471] | P[472] | P[473] | 
                    P[474] | P[475] | P[476] | P[477] | P[478] | P[479] | 
                    P[480] | P[481] | P[482] | P[483] | P[484] | P[485] | 
                    P[486] | P[487] | P[488] | P[489] | P[490] | P[491] | 
                    P[492] | P[493] | P[494] | P[495] | P[496] | P[497] | 
                    P[498] | P[499] | P[500] | P[501] | P[502] | P[503] | 
                    P[504] | P[505] | P[506] | P[507] | P[508] | P[509] | 
                    P[510] | P[511];
        Q[12] <= #1 P[  4] | P[  6] | P[ 13] | P[ 15] | P[ 17] | P[ 21] | 
                    P[ 23] | P[ 26] | P[ 28] | P[ 30] | P[ 34] | P[ 36] | 
                    P[ 38] | P[ 48] | P[ 50] | P[ 52] | P[ 54] | P[ 56] | 
                    P[ 58] | P[ 60] | P[ 62] | P[ 64] | P[ 66] | P[ 68] | 
                    P[ 70] | P[ 72] | P[ 74] | P[ 76] | P[ 78] | P[ 80] | 
                    P[ 82] | P[ 85] | P[ 87] | P[ 90] | P[ 92] | P[ 95] | 
                    P[ 97] | P[100] | P[102] | P[105] | P[107] | P[110] | 
                    P[112] | P[116] | P[117] | P[123] | P[125] | P[130] | 
                    P[134] | P[136] | P[138] | P[140] | P[142] | P[144] | 
                    P[150] | P[153] | P[159] | P[161] | P[166] | P[167] | 
                    P[170] | P[172] | P[174] | P[176] | P[186] | P[188] | 
                    P[189] | P[210] | P[215] | P[219];
        Q[13] <= #1 P[ 64] | P[ 82] | P[ 97] | P[112] | P[208];
        Q[14] <= #1 P[ 28] | P[ 30] | P[ 54] | P[ 56] | P[ 58] | P[ 72] | 
                    P[ 74] | P[ 76] | P[ 90] | P[ 92] | P[105] | P[107] | 
                    P[116] | P[123] | P[207] | P[210];
        Q[15] <= #1 P[  5] | P[ 14] | P[ 22] | P[ 29] | P[ 31] | P[ 32] | 
                    P[ 35] | P[ 37] | P[ 49] | P[ 51] | P[ 53] | P[ 55] | 
                    P[ 57] | P[ 59] | P[ 61] | P[ 63] | P[ 65] | P[ 67] | 
                    P[ 69] | P[ 71] | P[ 73] | P[ 75] | P[ 77] | P[ 79] | 
                    P[ 81] | P[ 83] | P[ 86] | P[ 88] | P[ 91] | P[ 93] | 
                    P[ 96] | P[ 98] | P[101] | P[103] | P[106] | P[108] | 
                    P[111] | P[113] | P[118] | P[119] | P[120] | P[121] | 
                    P[126] | P[127] | P[128] | P[129] | P[131] | P[132] | 
                    P[133] | P[135] | P[137] | P[139] | P[141] | P[162] | 
                    P[163] | P[164] | P[168] | P[171] | P[175] | P[178] | 
                    P[181] | P[182] | P[187] | P[192] | P[203] | P[204] | 
                    P[205] | P[206] | P[211] | P[212] | P[213] | P[214] | 
                    P[216] | P[217] | P[218] | P[220];
        Q[16] <= #1 P[184] | P[185] | P[194] | P[195] | P[196] | P[197] | 
                    P[198] | P[199] | P[200] | P[201] | P[202] | P[435];
        Q[17] <= #1 P[  1] | P[  2] | P[  3] | P[  9] | P[ 10] | P[ 11] | 
                    P[ 12] | P[ 19] | P[ 20] | P[ 24] | P[ 25] | P[ 40] | 
                    P[ 43] | P[ 44] | P[ 46] | P[ 47] | P[115] | P[151] | 
                    P[152] | P[154] | P[155] | P[157] | P[158] | P[165] | 
                    P[169] | P[177] | P[179] | P[180] | P[183] | P[190] | 
                    P[191] | P[193] | P[260] | P[262] | P[384] | P[386] | 
                    P[388] | P[390] | P[421] | P[423] | P[429] | P[431] | 
                    P[436] | P[438] | P[439];
        Q[18] <= #1 P[  8] | P[ 16] | P[ 17] | P[ 18] | P[ 27] | P[ 33] | 
                    P[ 39] | P[ 41] | P[ 42] | P[ 45] | P[ 84] | P[ 89] | 
                    P[ 94] | P[ 99] | P[104] | P[109] | P[114] | P[122] | 
                    P[124] | P[143] | P[144] | P[145] | P[146] | P[147] | 
                    P[148] | P[149] | P[150] | P[153] | P[156] | P[160] | 
                    P[173] | P[209] | P[256] | P[257] | P[258] | P[259] | 
                    P[261] | P[263] | P[264] | P[265] | P[266] | P[267] | 
                    P[268] | P[269] | P[270] | P[271] | P[272] | P[273] | 
                    P[274] | P[275] | P[276] | P[277] | P[278] | P[279] | 
                    P[280] | P[281] | P[282] | P[283] | P[284] | P[285] | 
                    P[286] | P[287] | P[288] | P[289] | P[290] | P[291] | 
                    P[292] | P[293] | P[294] | P[295] | P[296] | P[297] | 
                    P[298] | P[299] | P[300] | P[301] | P[302] | P[303] | 
                    P[304] | P[305] | P[306] | P[307] | P[308] | P[309] | 
                    P[310] | P[311] | P[312] | P[313] | P[314] | P[315] | 
                    P[316] | P[317] | P[318] | P[319] | P[320] | P[321] | 
                    P[322] | P[323] | P[324] | P[325] | P[326] | P[327] | 
                    P[328] | P[329] | P[330] | P[331] | P[332] | P[333] | 
                    P[334] | P[335] | P[336] | P[337] | P[338] | P[339] | 
                    P[340] | P[341] | P[342] | P[343] | P[344] | P[345] | 
                    P[346] | P[347] | P[348] | P[349] | P[350] | P[351] | 
                    P[352] | P[353] | P[354] | P[355] | P[356] | P[357] | 
                    P[358] | P[359] | P[360] | P[361] | P[362] | P[363] | 
                    P[364] | P[365] | P[366] | P[367] | P[368] | P[369] | 
                    P[370] | P[371] | P[372] | P[373] | P[374] | P[375] | 
                    P[376] | P[377] | P[378] | P[379] | P[380] | P[381] | 
                    P[382] | P[383] | P[385] | P[387] | P[389] | P[391] | 
                    P[392] | P[393] | P[394] | P[395] | P[396] | P[397] | 
                    P[398] | P[399] | P[400] | P[401] | P[402] | P[403] | 
                    P[404] | P[405] | P[406] | P[407] | P[408] | P[409] | 
                    P[410] | P[411] | P[412] | P[413] | P[414] | P[415] | 
                    P[416] | P[417] | P[418] | P[419] | P[420] | P[422] | 
                    P[424] | P[425] | P[426] | P[427] | P[428] | P[430] | 
                    P[432] | P[433] | P[434] | P[437] | P[440] | P[441] | 
                    P[442] | P[443] | P[444] | P[445] | P[446] | P[447] | 
                    P[448] | P[449] | P[450] | P[451] | P[452] | P[453] | 
                    P[454] | P[455] | P[456] | P[457] | P[458] | P[459] | 
                    P[460] | P[461] | P[462] | P[463] | P[464] | P[465] | 
                    P[466] | P[467] | P[468] | P[469] | P[470] | P[471] | 
                    P[472] | P[473] | P[474] | P[475] | P[476] | P[477] | 
                    P[478] | P[479] | P[480] | P[481] | P[482] | P[483] | 
                    P[484] | P[485] | P[486] | P[487] | P[488] | P[489] | 
                    P[490] | P[491] | P[492] | P[493] | P[494] | P[495] | 
                    P[496] | P[497] | P[498] | P[499] | P[500] | P[501] | 
                    P[502] | P[503] | P[504] | P[505] | P[506] | P[507] | 
                    P[508] | P[509] | P[510] | P[511];
        Q[19] <= #1 P[  6] | P[  8] | P[ 13] | P[ 15] | P[ 16] | P[ 17] | 
                    P[ 18] | P[ 23] | P[ 26] | P[ 27] | P[ 33] | P[ 38] | 
                    P[ 39] | P[ 41] | P[ 42] | P[ 45] | P[ 84] | P[ 89] | 
                    P[ 94] | P[ 99] | P[104] | P[109] | P[114] | P[122] | 
                    P[124] | P[143] | P[144] | P[145] | P[146] | P[147] | 
                    P[148] | P[149] | P[153] | P[156] | P[160] | P[173] | 
                    P[188] | P[189] | P[209] | P[256] | P[257] | P[258] | 
                    P[259] | P[261] | P[263] | P[264] | P[265] | P[266] | 
                    P[267] | P[268] | P[269] | P[270] | P[271] | P[272] | 
                    P[273] | P[274] | P[275] | P[276] | P[277] | P[278] | 
                    P[279] | P[280] | P[281] | P[282] | P[283] | P[284] | 
                    P[285] | P[286] | P[287] | P[288] | P[289] | P[290] | 
                    P[291] | P[292] | P[293] | P[294] | P[295] | P[296] | 
                    P[297] | P[298] | P[299] | P[300] | P[301] | P[302] | 
                    P[303] | P[304] | P[305] | P[306] | P[307] | P[308] | 
                    P[309] | P[310] | P[311] | P[312] | P[313] | P[314] | 
                    P[315] | P[316] | P[317] | P[318] | P[319] | P[320] | 
                    P[321] | P[322] | P[323] | P[324] | P[325] | P[326] | 
                    P[327] | P[328] | P[329] | P[330] | P[331] | P[332] | 
                    P[333] | P[334] | P[335] | P[336] | P[337] | P[338] | 
                    P[339] | P[340] | P[341] | P[342] | P[343] | P[344] | 
                    P[345] | P[346] | P[347] | P[348] | P[349] | P[350] | 
                    P[351] | P[352] | P[353] | P[354] | P[355] | P[356] | 
                    P[357] | P[358] | P[359] | P[360] | P[361] | P[362] | 
                    P[363] | P[364] | P[365] | P[366] | P[367] | P[368] | 
                    P[369] | P[370] | P[371] | P[372] | P[373] | P[374] | 
                    P[375] | P[376] | P[377] | P[378] | P[379] | P[380] | 
                    P[381] | P[382] | P[383] | P[385] | P[387] | P[389] | 
                    P[391] | P[392] | P[393] | P[394] | P[395] | P[396] | 
                    P[397] | P[398] | P[399] | P[400] | P[401] | P[402] | 
                    P[403] | P[404] | P[405] | P[406] | P[407] | P[408] | 
                    P[409] | P[410] | P[411] | P[412] | P[413] | P[414] | 
                    P[415] | P[416] | P[417] | P[418] | P[419] | P[420] | 
                    P[422] | P[424] | P[425] | P[426] | P[427] | P[428] | 
                    P[430] | P[432] | P[433] | P[434] | P[437] | P[440] | 
                    P[441] | P[442] | P[443] | P[444] | P[445] | P[446] | 
                    P[447] | P[448] | P[449] | P[450] | P[451] | P[452] | 
                    P[453] | P[454] | P[455] | P[456] | P[457] | P[458] | 
                    P[459] | P[460] | P[461] | P[462] | P[463] | P[464] | 
                    P[465] | P[466] | P[467] | P[468] | P[469] | P[470] | 
                    P[471] | P[472] | P[473] | P[474] | P[475] | P[476] | 
                    P[477] | P[478] | P[479] | P[480] | P[481] | P[482] | 
                    P[483] | P[484] | P[485] | P[486] | P[487] | P[488] | 
                    P[489] | P[490] | P[491] | P[492] | P[493] | P[494] | 
                    P[495] | P[496] | P[497] | P[498] | P[499] | P[500] | 
                    P[501] | P[502] | P[503] | P[504] | P[505] | P[506] | 
                    P[507] | P[508] | P[509] | P[510] | P[511];
        Q[20] <= #1 P[  1] | P[  2] | P[  3] | P[  9] | P[ 10] | P[ 11] | 
                    P[ 12] | P[ 19] | P[ 20] | P[ 24] | P[ 25] | P[ 40] | 
                    P[ 43] | P[ 44] | P[ 46] | P[ 47] | P[ 48] | P[ 49] | 
                    P[ 50] | P[ 51] | P[ 52] | P[ 53] | P[ 54] | P[ 55] | 
                    P[ 56] | P[ 57] | P[ 58] | P[ 59] | P[ 60] | P[ 61] | 
                    P[ 62] | P[ 63] | P[ 64] | P[ 65] | P[ 66] | P[ 67] | 
                    P[ 68] | P[ 69] | P[ 70] | P[ 71] | P[ 72] | P[ 73] | 
                    P[ 74] | P[ 75] | P[ 76] | P[ 77] | P[ 78] | P[ 79] | 
                    P[ 80] | P[ 81] | P[ 82] | P[ 83] | P[115] | P[116] | 
                    P[117] | P[118] | P[119] | P[120] | P[136] | P[137] | 
                    P[140] | P[141] | P[151] | P[152] | P[154] | P[155] | 
                    P[157] | P[158] | P[159] | P[162] | P[163] | P[164] | 
                    P[165] | P[169] | P[170] | P[171] | P[172] | P[177] | 
                    P[179] | P[180] | P[183] | P[190] | P[191] | P[193] | 
                    P[202] | P[203] | P[204] | P[205] | P[210] | P[211] | 
                    P[212] | P[213] | P[260] | P[262] | P[384] | P[386] | 
                    P[388] | P[390] | P[421] | P[423] | P[429] | P[431] | 
                    P[436] | P[438] | P[439];
        Q[21] <= #1 P[ 52] | P[ 58] | P[ 64] | P[ 70] | P[ 76] | P[ 82] | 
                    P[ 87] | P[ 92] | P[ 97] | P[102] | P[107] | P[112] | 
                    P[132] | P[183] | P[196] | P[200] | P[217] | P[388] | 
                    P[421] | P[429] | P[439];
        Q[22] <= #1 P[132] | P[217];
        Q[23] <= #1 P[ 48] | P[ 50] | P[ 52] | P[ 60] | P[ 62] | P[ 66] | 
                    P[ 68] | P[ 70] | P[ 78] | P[ 80] | P[ 85] | P[ 87] | 
                    P[ 95] | P[100] | P[102] | P[110] | P[116] | P[117] | 
                    P[125] | P[136] | P[140];
        Q[24] <= #1 P[  0] | P[  1] | P[  3] | P[  5] | P[  9] | P[ 10] | 
                    P[ 11] | P[ 13] | P[ 15] | P[ 17] | P[ 19] | P[ 20] | 
                    P[ 21] | P[ 23] | P[ 25] | P[ 35] | P[ 37] | P[ 40] | 
                    P[ 41] | P[ 43] | P[ 46] | P[ 47] | P[ 49] | P[ 51] | 
                    P[ 55] | P[ 57] | P[ 61] | P[ 63] | P[ 84] | P[ 85] | 
                    P[ 91] | P[ 94] | P[ 95] | P[101] | P[104] | P[105] | 
                    P[111] | P[131] | P[136] | P[137] | P[140] | P[141] | 
                    P[143] | P[145] | P[147] | P[149] | P[151] | P[153] | 
                    P[157] | P[162] | P[164] | P[166] | P[167] | P[169] | 
                    P[172] | P[175] | P[176] | P[177] | P[179] | P[181] | 
                    P[183] | P[187] | P[189] | P[193] | P[195] | P[202] | 
                    P[207] | P[208] | P[209] | P[210] | P[211] | P[212] | 
                    P[213] | P[215] | P[217] | P[219] | P[262] | P[266] | 
                    P[268] | P[270] | P[298] | P[300] | P[320] | P[321] | 
                    P[325] | P[333] | P[352] | P[354] | P[356] | P[358] | 
                    P[364] | P[366] | P[385] | P[387] | P[388] | P[389] | 
                    P[391] | P[393] | P[395] | P[397] | P[399] | P[400] | 
                    P[402] | P[404] | P[406] | P[408] | P[409] | P[410] | 
                    P[412] | P[414] | P[417] | P[419] | P[421] | P[425] | 
                    P[427] | P[429] | P[433] | P[435] | P[437] | P[438] | 
                    P[439] | P[441] | P[443] | P[445] | P[447] | P[451] | 
                    P[453] | P[454] | P[455] | P[456] | P[457] | P[459] | 
                    P[463] | P[465] | P[467] | P[469] | P[471] | P[472] | 
                    P[475] | P[477] | P[479] | P[488];
        Q[25] <= #1 P[  2] | P[  3] | P[  6] | P[  9] | P[ 10] | P[ 11] | 
                    P[ 14] | P[ 15] | P[ 18] | P[ 19] | P[ 22] | P[ 23] | 
                    P[ 26] | P[ 30] | P[ 31] | P[ 33] | P[ 34] | P[ 35] | 
                    P[ 38] | P[ 40] | P[ 41] | P[ 43] | P[ 44] | P[ 46] | 
                    P[ 50] | P[ 51] | P[ 54] | P[ 57] | P[ 61] | P[ 62] | 
                    P[ 66] | P[ 69] | P[ 74] | P[ 75] | P[ 78] | P[ 79] | 
                    P[ 86] | P[ 89] | P[ 90] | P[ 91] | P[ 94] | P[ 95] | 
                    P[106] | P[109] | P[110] | P[111] | P[114] | P[115] | 
                    P[116] | P[117] | P[118] | P[119] | P[121] | P[122] | 
                    P[123] | P[125] | P[126] | P[127] | P[129] | P[130] | 
                    P[131] | P[133] | P[134] | P[135] | P[138] | P[139] | 
                    P[142] | P[143] | P[148] | P[150] | P[151] | P[154] | 
                    P[159] | P[161] | P[162] | P[163] | P[167] | P[170] | 
                    P[173] | P[174] | P[179] | P[183] | P[185] | P[186] | 
                    P[193] | P[194] | P[195] | P[198] | P[199] | P[202] | 
                    P[203] | P[204] | P[206] | P[207] | P[208] | P[210] | 
                    P[211] | P[212] | P[215] | P[219] | P[256] | P[258] | 
                    P[266] | P[268] | P[270] | P[272] | P[274] | P[276] | 
                    P[278] | P[281] | P[282] | P[284] | P[286] | P[290] | 
                    P[294] | P[298] | P[300] | P[304] | P[305] | P[306] | 
                    P[307] | P[308] | P[309] | P[310] | P[311] | P[312] | 
                    P[313] | P[314] | P[315] | P[316] | P[317] | P[318] | 
                    P[319] | P[322] | P[324] | P[325] | P[327] | P[329] | 
                    P[330] | P[332] | P[333] | P[334] | P[336] | P[338] | 
                    P[340] | P[342] | P[345] | P[346] | P[348] | P[350] | 
                    P[362] | P[363] | P[387] | P[390] | P[391] | P[394] | 
                    P[395] | P[398] | P[399] | P[400] | P[401] | P[402] | 
                    P[403] | P[404] | P[405] | P[406] | P[407] | P[408] | 
                    P[410] | P[411] | P[412] | P[413] | P[414] | P[415] | 
                    P[418] | P[419] | P[422] | P[423] | P[426] | P[427] | 
                    P[430] | P[431] | P[434] | P[436] | P[438] | P[439] | 
                    P[442] | P[443] | P[446] | P[447] | P[455] | P[456] | 
                    P[457] | P[472] | P[481] | P[483] | P[485] | P[487] | 
                    P[488] | P[491] | P[493] | P[495];
        Q[26] <= #1 P[  4] | P[  5] | P[  6] | P[ 12] | P[ 13] | P[ 14] | 
                    P[ 15] | P[ 20] | P[ 21] | P[ 22] | P[ 23] | P[ 27] | 
                    P[ 28] | P[ 29] | P[ 30] | P[ 31] | P[ 32] | P[ 36] | 
                    P[ 37] | P[ 38] | P[ 41] | P[ 47] | P[ 49] | P[ 51] | 
                    P[ 54] | P[ 55] | P[ 57] | P[ 60] | P[ 61] | P[ 62] | 
                    P[ 67] | P[ 68] | P[ 69] | P[ 73] | P[ 75] | P[ 78] | 
                    P[ 79] | P[ 84] | P[ 85] | P[ 86] | P[ 91] | P[ 94] | 
                    P[ 95] | P[ 99] | P[100] | P[101] | P[106] | P[109] | 
                    P[110] | P[111] | P[116] | P[117] | P[119] | P[120] | 
                    P[123] | P[124] | P[125] | P[127] | P[128] | P[132] | 
                    P[134] | P[140] | P[141] | P[142] | P[143] | P[149] | 
                    P[151] | P[156] | P[157] | P[162] | P[163] | P[166] | 
                    P[167] | P[169] | P[173] | P[174] | P[180] | P[181] | 
                    P[183] | P[187] | P[188] | P[189] | P[195] | P[198] | 
                    P[199] | P[204] | P[205] | P[207] | P[208] | P[211] | 
                    P[215] | P[266] | P[268] | P[270] | P[272] | P[273] | 
                    P[274] | P[275] | P[276] | P[277] | P[278] | P[279] | 
                    P[281] | P[282] | P[283] | P[284] | P[285] | P[286] | 
                    P[287] | P[292] | P[294] | P[297] | P[298] | P[300] | 
                    P[302] | P[312] | P[320] | P[321] | P[325] | P[326] | 
                    P[328] | P[333] | P[335] | P[344] | P[352] | P[353] | 
                    P[354] | P[355] | P[356] | P[357] | P[358] | P[359] | 
                    P[360] | P[363] | P[364] | P[365] | P[366] | P[367] | 
                    P[388] | P[389] | P[391] | P[396] | P[397] | P[398] | 
                    P[399] | P[400] | P[401] | P[402] | P[403] | P[404] | 
                    P[405] | P[406] | P[407] | P[408] | P[409] | P[410] | 
                    P[411] | P[412] | P[413] | P[414] | P[415] | P[420] | 
                    P[421] | P[422] | P[428] | P[429] | P[430] | P[436] | 
                    P[437] | P[438] | P[439] | P[444] | P[445] | P[446] | 
                    P[447] | P[448] | P[449] | P[450] | P[453] | P[458] | 
                    P[460] | P[462] | P[463] | P[464] | P[466] | P[468] | 
                    P[470] | P[474] | P[476] | P[478] | P[480] | P[482] | 
                    P[484] | P[486] | P[490] | P[491] | P[492] | P[494] | 
                    P[496] | P[497] | P[498] | P[499] | P[500] | P[501] | 
                    P[502] | P[503] | P[504] | P[505] | P[506] | P[507] | 
                    P[508] | P[509] | P[510] | P[511];
        Q[27] <= #1 P[  8] | P[  9] | P[ 10] | P[ 11] | P[ 12] | P[ 13] | 
                    P[ 14] | P[ 15] | P[ 24] | P[ 25] | P[ 26] | P[ 27] | 
                    P[ 28] | P[ 30] | P[ 39] | P[ 40] | P[ 42] | P[ 43] | 
                    P[ 44] | P[ 45] | P[ 46] | P[ 47] | P[ 52] | P[ 53] | 
                    P[ 56] | P[ 58] | P[ 59] | P[ 60] | P[ 61] | P[ 62] | 
                    P[ 64] | P[ 65] | P[ 70] | P[ 71] | P[ 72] | P[ 74] | 
                    P[ 76] | P[ 77] | P[ 78] | P[ 79] | P[ 82] | P[ 83] | 
                    P[ 87] | P[ 88] | P[ 89] | P[ 90] | P[ 92] | P[ 93] | 
                    P[ 94] | P[ 95] | P[ 97] | P[ 98] | P[102] | P[103] | 
                    P[104] | P[105] | P[107] | P[108] | P[109] | P[110] | 
                    P[111] | P[112] | P[113] | P[115] | P[122] | P[123] | 
                    P[124] | P[125] | P[136] | P[137] | P[138] | P[140] | 
                    P[141] | P[142] | P[143] | P[146] | P[147] | P[150] | 
                    P[152] | P[153] | P[154] | P[155] | P[156] | P[157] | 
                    P[158] | P[164] | P[165] | P[168] | P[170] | P[173] | 
                    P[174] | P[178] | P[182] | P[184] | P[185] | P[186] | 
                    P[187] | P[188] | P[189] | P[190] | P[193] | P[196] | 
                    P[197] | P[200] | P[201] | P[202] | P[207] | P[208] | 
                    P[212] | P[213] | P[214] | P[216] | P[217] | P[218] | 
                    P[219] | P[220] | P[256] | P[260] | P[262] | P[273] | 
                    P[275] | P[277] | P[279] | P[280] | P[281] | P[283] | 
                    P[285] | P[287] | P[288] | P[296] | P[302] | P[305] | 
                    P[307] | P[309] | P[311] | P[313] | P[315] | P[317] | 
                    P[319] | P[323] | P[325] | P[327] | P[329] | P[331] | 
                    P[333] | P[335] | P[337] | P[339] | P[341] | P[343] | 
                    P[345] | P[347] | P[349] | P[351] | P[363] | P[368] | 
                    P[369] | P[370] | P[371] | P[372] | P[373] | P[374] | 
                    P[375] | P[376] | P[377] | P[378] | P[379] | P[380] | 
                    P[381] | P[382] | P[383] | P[384] | P[386] | P[388] | 
                    P[390] | P[392] | P[393] | P[394] | P[395] | P[396] | 
                    P[397] | P[398] | P[399] | P[401] | P[403] | P[405] | 
                    P[407] | P[409] | P[411] | P[413] | P[415] | P[421] | 
                    P[423] | P[424] | P[425] | P[426] | P[427] | P[428] | 
                    P[429] | P[430] | P[431] | P[435] | P[436] | P[438] | 
                    P[440] | P[441] | P[442] | P[443] | P[444] | P[445] | 
                    P[446] | P[447] | P[448] | P[449] | P[451] | P[455] | 
                    P[459] | P[463] | P[465] | P[467] | P[469] | P[471] | 
                    P[473] | P[475] | P[477] | P[479] | P[480] | P[481] | 
                    P[482] | P[483] | P[484] | P[485] | P[486] | P[487] | 
                    P[489] | P[491] | P[492] | P[493] | P[494] | P[495] | 
                    P[496] | P[497] | P[498] | P[499] | P[500] | P[501] | 
                    P[502] | P[503] | P[504] | P[505] | P[506] | P[507] | 
                    P[508] | P[509] | P[510] | P[511];
        Q[28] <= #1 P[ 16] | P[ 17] | P[ 18] | P[ 19] | P[ 20] | P[ 21] | 
                    P[ 22] | P[ 23] | P[ 24] | P[ 25] | P[ 26] | P[ 27] | 
                    P[ 28] | P[ 30] | P[ 48] | P[ 49] | P[ 50] | P[ 51] | 
                    P[ 54] | P[ 55] | P[ 56] | P[ 57] | P[ 60] | P[ 61] | 
                    P[ 62] | P[ 80] | P[ 81] | P[ 84] | P[ 85] | P[ 86] | 
                    P[ 89] | P[ 90] | P[ 91] | P[ 94] | P[ 95] | P[114] | 
                    P[116] | P[117] | P[121] | P[122] | P[123] | P[124] | 
                    P[125] | P[129] | P[133] | P[135] | P[139] | P[144] | 
                    P[145] | P[148] | P[149] | P[150] | P[151] | P[152] | 
                    P[153] | P[154] | P[156] | P[157] | P[171] | P[172] | 
                    P[175] | P[176] | P[177] | P[179] | P[180] | P[181] | 
                    P[183] | P[184] | P[185] | P[186] | P[187] | P[188] | 
                    P[189] | P[195] | P[206] | P[209] | P[210] | P[211] | 
                    P[212] | P[213] | P[215] | P[216] | P[217] | P[219] | 
                    P[257] | P[258] | P[259] | P[260] | P[261] | P[262] | 
                    P[263] | P[264] | P[265] | P[267] | P[269] | P[271] | 
                    P[272] | P[273] | P[274] | P[275] | P[276] | P[277] | 
                    P[278] | P[279] | P[282] | P[283] | P[284] | P[285] | 
                    P[286] | P[287] | P[289] | P[291] | P[293] | P[295] | 
                    P[299] | P[301] | P[302] | P[303] | P[320] | P[321] | 
                    P[322] | P[323] | P[324] | P[330] | P[331] | P[332] | 
                    P[333] | P[334] | P[336] | P[337] | P[338] | P[339] | 
                    P[340] | P[341] | P[342] | P[343] | P[346] | P[347] | 
                    P[348] | P[349] | P[350] | P[351] | P[352] | P[353] | 
                    P[354] | P[355] | P[356] | P[357] | P[358] | P[359] | 
                    P[361] | P[362] | P[363] | P[364] | P[365] | P[366] | 
                    P[367] | P[401] | P[403] | P[405] | P[407] | P[411] | 
                    P[413] | P[415] | P[432] | P[433] | P[434] | P[435] | 
                    P[436] | P[437] | P[438] | P[439] | P[440] | P[441] | 
                    P[442] | P[443] | P[444] | P[445] | P[446] | P[447] | 
                    P[448] | P[449] | P[450] | P[451] | P[453] | P[455] | 
                    P[458] | P[459] | P[460] | P[462] | P[464] | P[465] | 
                    P[466] | P[467] | P[468] | P[469] | P[470] | P[471] | 
                    P[474] | P[475] | P[476] | P[477] | P[478] | P[479] | 
                    P[480] | P[481] | P[482] | P[483] | P[484] | P[485] | 
                    P[486] | P[487] | P[490] | P[491] | P[492] | P[493] | 
                    P[494] | P[495];
        Q[29] <= #1 P[ 29] | P[ 31] | P[ 32] | P[ 33] | P[ 34] | P[ 35] | 
                    P[ 36] | P[ 37] | P[ 38] | P[ 41] | P[ 44] | P[ 47] | 
                    P[ 48] | P[ 50] | P[ 54] | P[ 56] | P[ 60] | P[ 62] | 
                    P[ 63] | P[ 67] | P[ 69] | P[ 73] | P[ 75] | P[ 79] | 
                    P[ 81] | P[ 96] | P[ 99] | P[100] | P[101] | P[104] | 
                    P[105] | P[106] | P[109] | P[110] | P[111] | P[114] | 
                    P[116] | P[117] | P[121] | P[122] | P[123] | P[124] | 
                    P[125] | P[129] | P[133] | P[135] | P[139] | P[159] | 
                    P[160] | P[161] | P[162] | P[163] | P[164] | P[166] | 
                    P[167] | P[168] | P[169] | P[170] | P[171] | P[172] | 
                    P[173] | P[174] | P[175] | P[176] | P[177] | P[179] | 
                    P[180] | P[181] | P[183] | P[184] | P[185] | P[186] | 
                    P[187] | P[188] | P[189] | P[199] | P[206] | P[266] | 
                    P[268] | P[270] | P[272] | P[273] | P[274] | P[275] | 
                    P[276] | P[277] | P[278] | P[279] | P[282] | P[283] | 
                    P[284] | P[285] | P[286] | P[287] | P[289] | P[290] | 
                    P[291] | P[292] | P[293] | P[294] | P[295] | P[296] | 
                    P[298] | P[299] | P[300] | P[301] | P[303] | P[320] | 
                    P[321] | P[322] | P[323] | P[330] | P[331] | P[332] | 
                    P[334] | P[335] | P[336] | P[337] | P[338] | P[339] | 
                    P[340] | P[341] | P[342] | P[343] | P[346] | P[347] | 
                    P[348] | P[349] | P[350] | P[351] | P[352] | P[353] | 
                    P[354] | P[355] | P[356] | P[357] | P[358] | P[359] | 
                    P[362] | P[363] | P[364] | P[365] | P[366] | P[367] | 
                    P[388] | P[390] | P[400] | P[402] | P[404] | P[406] | 
                    P[408] | P[409] | P[410] | P[412] | P[414] | P[416] | 
                    P[417] | P[418] | P[419] | P[420] | P[421] | P[422] | 
                    P[423] | P[424] | P[425] | P[426] | P[427] | P[428] | 
                    P[429] | P[430] | P[431] | P[432] | P[433] | P[434] | 
                    P[435] | P[436] | P[437] | P[438] | P[439] | P[440] | 
                    P[441] | P[442] | P[443] | P[444] | P[445] | P[446] | 
                    P[447] | P[448] | P[449] | P[452] | P[454] | P[456] | 
                    P[457] | P[461] | P[463] | P[472] | P[473] | P[480] | 
                    P[481] | P[482] | P[483] | P[484] | P[485] | P[486] | 
                    P[487] | P[488] | P[489] | P[492] | P[493] | P[494] | 
                    P[495];
        Q[30] <= #1 P[ 49] | P[ 51] | P[ 55] | P[ 57] | P[ 61] | P[ 63] | 
                    P[ 66] | P[ 67] | P[ 68] | P[ 69] | P[ 72] | P[ 73] | 
                    P[ 74] | P[ 75] | P[ 78] | P[ 79] | P[ 80] | P[ 81] | 
                    P[ 84] | P[ 85] | P[ 86] | P[ 89] | P[ 90] | P[ 91] | 
                    P[ 94] | P[ 95] | P[ 96] | P[ 99] | P[100] | P[101] | 
                    P[104] | P[105] | P[106] | P[109] | P[110] | P[111] | 
                    P[114] | P[116] | P[117] | P[121] | P[122] | P[123] | 
                    P[124] | P[125] | P[129] | P[133] | P[135] | P[139] | 
                    P[191] | P[192] | P[194] | P[195] | P[198] | P[199] | 
                    P[202] | P[206] | P[207] | P[208] | P[209] | P[210] | 
                    P[211] | P[212] | P[213] | P[215] | P[216] | P[217] | 
                    P[219] | P[280] | P[281] | P[297] | P[304] | P[305] | 
                    P[306] | P[307] | P[308] | P[309] | P[310] | P[311] | 
                    P[312] | P[313] | P[314] | P[315] | P[316] | P[317] | 
                    P[318] | P[319] | P[320] | P[321] | P[324] | P[325] | 
                    P[326] | P[327] | P[328] | P[329] | P[344] | P[345] | 
                    P[352] | P[353] | P[354] | P[355] | P[356] | P[357] | 
                    P[358] | P[359] | P[360] | P[361] | P[364] | P[365] | 
                    P[366] | P[367] | P[401] | P[403] | P[405] | P[407] | 
                    P[409] | P[411] | P[413] | P[415] | P[448] | P[449] | 
                    P[450] | P[451] | P[456] | P[457] | P[458] | P[459] | 
                    P[460] | P[462] | P[464] | P[465] | P[466] | P[467] | 
                    P[468] | P[469] | P[470] | P[471] | P[472] | P[473] | 
                    P[474] | P[475] | P[476] | P[477] | P[478] | P[479] | 
                    P[480] | P[481] | P[482] | P[483] | P[484] | P[485] | 
                    P[486] | P[487] | P[488] | P[489] | P[490] | P[491] | 
                    P[492] | P[493] | P[494] | P[495];
        Q[31] <= #1 P[118] | P[119] | P[120] | P[126] | P[127] | P[128] | 
                    P[130] | P[131] | P[132] | P[134] | P[136] | P[137] | 
                    P[138] | P[140] | P[141] | P[142] | P[143] | P[144] | 
                    P[145] | P[148] | P[149] | P[150] | P[151] | P[152] | 
                    P[153] | P[154] | P[156] | P[157] | P[159] | P[160] | 
                    P[161] | P[162] | P[163] | P[164] | P[166] | P[167] | 
                    P[168] | P[169] | P[170] | P[171] | P[172] | P[173] | 
                    P[174] | P[175] | P[176] | P[177] | P[179] | P[180] | 
                    P[181] | P[183] | P[184] | P[185] | P[186] | P[187] | 
                    P[188] | P[189] | P[191] | P[192] | P[194] | P[198] | 
                    P[202] | P[203] | P[204] | P[205] | P[207] | P[208] | 
                    P[209] | P[210] | P[211] | P[212] | P[213] | P[215] | 
                    P[216] | P[217] | P[219] | P[302] | P[304] | P[305] | 
                    P[306] | P[307] | P[308] | P[309] | P[310] | P[311] | 
                    P[312] | P[313] | P[314] | P[315] | P[316] | P[317] | 
                    P[318] | P[319] | P[324] | P[325] | P[333] | P[335] | 
                    P[368] | P[369] | P[370] | P[371] | P[372] | P[373] | 
                    P[374] | P[375] | P[376] | P[377] | P[378] | P[379] | 
                    P[380] | P[381] | P[382] | P[383] | P[385] | P[387] | 
                    P[389] | P[391] | P[392] | P[393] | P[394] | P[395] | 
                    P[396] | P[397] | P[398] | P[399] | P[416] | P[417] | 
                    P[418] | P[419] | P[420] | P[422] | P[424] | P[425] | 
                    P[426] | P[427] | P[428] | P[430] | P[432] | P[433] | 
                    P[434] | P[435] | P[436] | P[437] | P[438] | P[439] | 
                    P[440] | P[441] | P[442] | P[443] | P[444] | P[445] | 
                    P[446] | P[447] | P[453] | P[461] | P[463] | P[496] | 
                    P[497] | P[498] | P[499] | P[500] | P[501] | P[502] | 
                    P[503] | P[504] | P[505] | P[506] | P[507] | P[508] | 
                    P[509] | P[510] | P[511];
        Q[32] <= #1 P[  6] | P[  8] | P[ 15] | P[ 17] | P[ 23] | P[ 26] | 
                    P[ 38] | P[ 39] | P[ 41] | P[ 42] | P[ 44] | P[ 45] | 
                    P[ 47] | P[ 52] | P[ 53] | P[ 58] | P[ 59] | P[ 64] | 
                    P[ 65] | P[ 70] | P[ 71] | P[ 76] | P[ 77] | P[ 82] | 
                    P[ 83] | P[ 87] | P[ 88] | P[ 92] | P[ 93] | P[ 97] | 
                    P[ 98] | P[102] | P[103] | P[107] | P[108] | P[112] | 
                    P[113] | P[114] | P[116] | P[117] | P[121] | P[123] | 
                    P[125] | P[129] | P[133] | P[135] | P[139] | P[144] | 
                    P[146] | P[148] | P[153] | P[155] | P[158] | P[159] | 
                    P[161] | P[165] | P[178] | P[182] | P[188] | P[189] | 
                    P[190] | P[191] | P[192] | P[196] | P[197] | P[200] | 
                    P[201] | P[202] | P[206] | P[209] | P[210] | P[214] | 
                    P[218] | P[220] | P[257] | P[259] | P[261] | P[263] | 
                    P[264] | P[265] | P[267] | P[269] | P[271] | P[288] | 
                    P[290] | P[292] | P[294] | P[296] | P[384] | P[385] | 
                    P[386] | P[387] | P[389] | P[391] | P[392] | P[393] | 
                    P[394] | P[395] | P[396] | P[397] | P[398] | P[399] | 
                    P[416] | P[417] | P[418] | P[419] | P[420] | P[422] | 
                    P[424] | P[425] | P[426] | P[427] | P[428] | P[430] | 
                    P[432] | P[433] | P[434] | P[437] | P[440] | P[441] | 
                    P[442] | P[443] | P[444] | P[445] | P[446] | P[447];
        Q[33] <= #1 P[  0] | P[  1] | P[  2] | P[  3] | P[  4] | P[  5] | 
                    P[  9] | P[ 10] | P[ 11] | P[ 12] | P[ 13] | P[ 14] | 
                    P[ 16] | P[ 18] | P[ 19] | P[ 20] | P[ 21] | P[ 22] | 
                    P[ 24] | P[ 25] | P[ 27] | P[ 28] | P[ 30] | P[ 31] | 
                    P[ 32] | P[ 33] | P[ 34] | P[ 35] | P[ 36] | P[ 37] | 
                    P[ 40] | P[ 41] | P[ 43] | P[ 44] | P[ 46] | P[ 47] | 
                    P[ 48] | P[ 50] | P[ 52] | P[ 53] | P[ 54] | P[ 56] | 
                    P[ 58] | P[ 59] | P[ 60] | P[ 62] | P[ 64] | P[ 65] | 
                    P[ 66] | P[ 68] | P[ 70] | P[ 71] | P[ 72] | P[ 74] | 
                    P[ 76] | P[ 77] | P[ 78] | P[ 80] | P[ 82] | P[ 83] | 
                    P[ 84] | P[ 85] | P[ 86] | P[ 87] | P[ 88] | P[ 89] | 
                    P[ 90] | P[ 92] | P[ 93] | P[ 94] | P[ 95] | P[ 96] | 
                    P[ 97] | P[ 98] | P[ 99] | P[100] | P[101] | P[102] | 
                    P[103] | P[104] | P[105] | P[107] | P[108] | P[109] | 
                    P[110] | P[111] | P[112] | P[113] | P[115] | P[121] | 
                    P[122] | P[124] | P[129] | P[130] | P[131] | P[132] | 
                    P[133] | P[134] | P[135] | P[136] | P[137] | P[138] | 
                    P[139] | P[140] | P[141] | P[142] | P[143] | P[146] | 
                    P[147] | P[148] | P[149] | P[151] | P[152] | P[154] | 
                    P[155] | P[156] | P[157] | P[158] | P[160] | P[165] | 
                    P[167] | P[168] | P[170] | P[173] | P[174] | P[177] | 
                    P[178] | P[179] | P[180] | P[181] | P[182] | P[183] | 
                    P[184] | P[185] | P[186] | P[190] | P[191] | P[193] | 
                    P[194] | P[196] | P[197] | P[198] | P[200] | P[201] | 
                    P[206] | P[207] | P[214] | P[215] | P[216] | P[218] | 
                    P[219] | P[220] | P[257] | P[259] | P[261] | P[263] | 
                    P[264] | P[265] | P[267] | P[269] | P[271] | P[272] | 
                    P[273] | P[274] | P[275] | P[276] | P[277] | P[278] | 
                    P[279] | P[280] | P[281] | P[282] | P[283] | P[284] | 
                    P[285] | P[286] | P[287] | P[288] | P[289] | P[290] | 
                    P[291] | P[292] | P[293] | P[294] | P[295] | P[296] | 
                    P[299] | P[301] | P[303] | P[304] | P[306] | P[308] | 
                    P[310] | P[312] | P[314] | P[316] | P[318] | P[322] | 
                    P[323] | P[326] | P[327] | P[328] | P[329] | P[330] | 
                    P[331] | P[332] | P[333] | P[334] | P[335] | P[336] | 
                    P[337] | P[338] | P[339] | P[340] | P[341] | P[342] | 
                    P[343] | P[344] | P[345] | P[346] | P[347] | P[348] | 
                    P[349] | P[350] | P[351] | P[360] | P[361] | P[362] | 
                    P[363] | P[384] | P[385] | P[386] | P[387] | P[392] | 
                    P[393] | P[394] | P[395] | P[396] | P[397] | P[398] | 
                    P[399] | P[416] | P[417] | P[418] | P[419] | P[420] | 
                    P[422] | P[424] | P[425] | P[426] | P[427] | P[428] | 
                    P[430] | P[432] | P[433] | P[434] | P[437] | P[453];
        Q[34] <= #1 P[  0] | P[  6] | P[  8] | P[  9] | P[ 10] | P[ 15] | 
                    P[ 17] | P[ 20] | P[ 23] | P[ 26] | P[ 27] | P[ 29] | 
                    P[ 32] | P[ 33] | P[ 38] | P[ 39] | P[ 40] | P[ 42] | 
                    P[ 43] | P[ 45] | P[ 46] | P[ 49] | P[ 51] | P[ 55] | 
                    P[ 57] | P[ 61] | P[ 63] | P[ 67] | P[ 69] | P[ 73] | 
                    P[ 75] | P[ 79] | P[ 81] | P[ 84] | P[ 89] | P[ 91] | 
                    P[ 94] | P[ 99] | P[104] | P[106] | P[109] | P[114] | 
                    P[115] | P[116] | P[117] | P[118] | P[119] | P[120] | 
                    P[123] | P[125] | P[126] | P[127] | P[128] | P[136] | 
                    P[140] | P[144] | P[145] | P[150] | P[153] | P[159] | 
                    P[161] | P[162] | P[163] | P[164] | P[166] | P[169] | 
                    P[171] | P[172] | P[173] | P[175] | P[176] | P[185] | 
                    P[187] | P[188] | P[189] | P[192] | P[193] | P[195] | 
                    P[199] | P[202] | P[203] | P[204] | P[205] | P[209] | 
                    P[210] | P[211] | P[212] | P[213] | P[217] | P[256] | 
                    P[257] | P[258] | P[259] | P[260] | P[261] | P[262] | 
                    P[263] | P[264] | P[265] | P[266] | P[267] | P[268] | 
                    P[269] | P[270] | P[271] | P[272] | P[273] | P[274] | 
                    P[275] | P[276] | P[277] | P[278] | P[279] | P[280] | 
                    P[281] | P[282] | P[283] | P[284] | P[285] | P[286] | 
                    P[287] | P[289] | P[290] | P[291] | P[292] | P[293] | 
                    P[294] | P[295] | P[296] | P[297] | P[298] | P[299] | 
                    P[300] | P[301] | P[302] | P[303] | P[304] | P[305] | 
                    P[306] | P[307] | P[308] | P[309] | P[310] | P[311] | 
                    P[312] | P[313] | P[314] | P[315] | P[316] | P[317] | 
                    P[318] | P[319] | P[320] | P[321] | P[322] | P[323] | 
                    P[324] | P[325] | P[326] | P[327] | P[328] | P[329] | 
                    P[330] | P[331] | P[332] | P[333] | P[334] | P[335] | 
                    P[336] | P[337] | P[338] | P[339] | P[340] | P[341] | 
                    P[342] | P[343] | P[344] | P[345] | P[346] | P[347] | 
                    P[348] | P[349] | P[350] | P[351] | P[352] | P[353] | 
                    P[354] | P[355] | P[356] | P[357] | P[358] | P[359] | 
                    P[360] | P[361] | P[362] | P[363] | P[364] | P[365] | 
                    P[366] | P[367] | P[368] | P[369] | P[370] | P[371] | 
                    P[372] | P[373] | P[374] | P[375] | P[376] | P[377] | 
                    P[378] | P[379] | P[380] | P[381] | P[382] | P[383] | 
                    P[385] | P[387] | P[388] | P[389] | P[390] | P[391] | 
                    P[392] | P[393] | P[394] | P[395] | P[396] | P[397] | 
                    P[398] | P[399] | P[400] | P[401] | P[402] | P[403] | 
                    P[404] | P[405] | P[406] | P[407] | P[408] | P[409] | 
                    P[410] | P[411] | P[412] | P[413] | P[414] | P[415] | 
                    P[416] | P[417] | P[418] | P[419] | P[420] | P[421] | 
                    P[422] | P[423] | P[424] | P[425] | P[426] | P[427] | 
                    P[428] | P[429] | P[430] | P[431] | P[432] | P[433] | 
                    P[434] | P[435] | P[436] | P[437] | P[438] | P[439] | 
                    P[440] | P[441] | P[442] | P[443] | P[444] | P[445] | 
                    P[446] | P[447] | P[448] | P[449] | P[450] | P[451] | 
                    P[452] | P[453] | P[454] | P[455] | P[456] | P[457] | 
                    P[458] | P[459] | P[460] | P[461] | P[462] | P[463] | 
                    P[464] | P[465] | P[466] | P[467] | P[468] | P[469] | 
                    P[470] | P[471] | P[472] | P[473] | P[474] | P[475] | 
                    P[476] | P[477] | P[478] | P[479] | P[480] | P[481] | 
                    P[482] | P[483] | P[484] | P[485] | P[486] | P[487] | 
                    P[488] | P[489] | P[490] | P[491] | P[492] | P[493] | 
                    P[494] | P[495] | P[496] | P[497] | P[498] | P[499] | 
                    P[500] | P[501] | P[502] | P[503] | P[504] | P[505] | 
                    P[506] | P[507] | P[508] | P[509] | P[510] | P[511];
        Q[35] <= #1 P[ 20] | P[ 27] | P[ 32] | P[ 33] | P[ 84] | P[ 89] | 
                    P[ 94] | P[ 99] | P[104] | P[109] | P[116] | P[117] | 
                    P[123] | P[125] | P[136] | P[140] | P[146] | P[147] | 
                    P[159] | P[161] | P[172] | P[173] | P[175] | P[176] | 
                    P[185] | P[202] | P[208] | P[210] | P[257] | P[259] | 
                    P[261] | P[263] | P[264] | P[265] | P[266] | P[267] | 
                    P[268] | P[269] | P[270] | P[271] | P[272] | P[273] | 
                    P[274] | P[275] | P[276] | P[277] | P[278] | P[279] | 
                    P[280] | P[281] | P[282] | P[283] | P[284] | P[285] | 
                    P[286] | P[287] | P[289] | P[291] | P[293] | P[295] | 
                    P[298] | P[299] | P[300] | P[301] | P[302] | P[303] | 
                    P[304] | P[306] | P[308] | P[310] | P[312] | P[314] | 
                    P[316] | P[318] | P[322] | P[323] | P[326] | P[327] | 
                    P[328] | P[329] | P[330] | P[331] | P[332] | P[333] | 
                    P[334] | P[335] | P[336] | P[337] | P[338] | P[339] | 
                    P[340] | P[341] | P[342] | P[343] | P[344] | P[345] | 
                    P[346] | P[347] | P[348] | P[349] | P[350] | P[351] | 
                    P[360] | P[361] | P[362] | P[363] | P[388] | P[390] | 
                    P[400] | P[402] | P[404] | P[406] | P[408] | P[410] | 
                    P[412] | P[414] | P[421] | P[423] | P[429] | P[431] | 
                    P[453];
    end
end

endmodule
